-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity dup2_0CLK_e4095020 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dup2_0CLK_e4095020;
architecture arch of dup2_0CLK_e4095020 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2790_c6_3167]
signal BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2790_c2_d3ad]
signal t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2790_c2_d3ad]
signal t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2790_c2_d3ad]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2790_c2_d3ad]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2790_c2_d3ad]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2790_c2_d3ad]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2790_c2_d3ad]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2790_c2_d3ad]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2790_c2_d3ad]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2790_c2_d3ad]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2790_c2_d3ad]
signal result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2803_c11_0552]
signal BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2803_c7_97e8]
signal t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2803_c7_97e8]
signal t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2803_c7_97e8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2803_c7_97e8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2803_c7_97e8]
signal result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2803_c7_97e8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2803_c7_97e8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2806_c11_aefa]
signal BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2806_c7_c4ed]
signal t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2806_c7_c4ed]
signal t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2806_c7_c4ed]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2806_c7_c4ed]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2806_c7_c4ed]
signal result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2806_c7_c4ed]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2806_c7_c4ed]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2808_c30_ca18]
signal sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2813_c11_8072]
signal BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2813_c7_63d9]
signal t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2813_c7_63d9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2813_c7_63d9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2813_c7_63d9]
signal result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2813_c7_63d9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2819_c11_f6eb]
signal BIN_OP_EQ_uxn_opcodes_h_l2819_c11_f6eb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2819_c11_f6eb_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2819_c11_f6eb_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2819_c7_5956]
signal result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2819_c7_5956]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2819_c7_5956]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2823_c11_72b9]
signal BIN_OP_EQ_uxn_opcodes_h_l2823_c11_72b9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2823_c11_72b9_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2823_c11_72b9_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2823_c7_c9e1]
signal result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2823_c7_c9e1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2823_c7_c9e1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8b52( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_opc_done := ref_toks_6;
      base.is_ram_write := ref_toks_7;
      base.is_vram_write := ref_toks_8;
      base.u8_value := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167
BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_left,
BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_right,
BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad
t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond,
t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue,
t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse,
t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad
t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond,
t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue,
t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse,
t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad
result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad
result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad
result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad
result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad
result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad
result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad
result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond,
result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552
BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_left,
BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_right,
BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8
t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_cond,
t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue,
t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse,
t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8
t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_cond,
t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue,
t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse,
t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8
result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8
result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8
result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_cond,
result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8
result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa
BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_left,
BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_right,
BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed
t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond,
t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue,
t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse,
t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed
t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond,
t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue,
t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse,
t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed
result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed
result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed
result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond,
result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed
result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18
sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_ins,
sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_x,
sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_y,
sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072
BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072_left,
BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072_right,
BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9
t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_cond,
t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue,
t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse,
t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9
result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9
result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_cond,
result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9
result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2819_c11_f6eb
BIN_OP_EQ_uxn_opcodes_h_l2819_c11_f6eb : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2819_c11_f6eb_left,
BIN_OP_EQ_uxn_opcodes_h_l2819_c11_f6eb_right,
BIN_OP_EQ_uxn_opcodes_h_l2819_c11_f6eb_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956
result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_cond,
result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956
result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2823_c11_72b9
BIN_OP_EQ_uxn_opcodes_h_l2823_c11_72b9 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2823_c11_72b9_left,
BIN_OP_EQ_uxn_opcodes_h_l2823_c11_72b9_right,
BIN_OP_EQ_uxn_opcodes_h_l2823_c11_72b9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1
result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_cond,
result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1
result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_return_output,
 t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output,
 t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_return_output,
 t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output,
 t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_return_output,
 t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output,
 t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output,
 sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072_return_output,
 t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2819_c11_f6eb_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2823_c11_72b9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2795_c3_4584 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2790_c2_d3ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2790_c2_d3ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2800_c3_1b36 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2790_c2_d3ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2790_c2_d3ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2804_c3_3a05 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2810_c3_5238 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2816_c3_7af6 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2815_c3_bc78 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2819_c11_f6eb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2819_c11_f6eb_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2819_c11_f6eb_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2820_c3_47e7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_72b9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_72b9_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_72b9_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2824_c3_2597 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2823_c7_c9e1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2803_l2823_l2790_DUPLICATE_c360_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2803_l2813_DUPLICATE_db7f_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2803_l2806_DUPLICATE_f768_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2819_l2813_l2806_l2803_l2823_DUPLICATE_1f5c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2829_l2786_DUPLICATE_f68a_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2819_c11_f6eb_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2810_c3_5238 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2810_c3_5238;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072_right := to_unsigned(3, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2815_c3_bc78 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2815_c3_bc78;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_right := to_unsigned(2, 2);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2800_c3_1b36 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2800_c3_1b36;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_right := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2824_c3_2597 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2824_c3_2597;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2804_c3_3a05 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2804_c3_3a05;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_iftrue := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2816_c3_7af6 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2816_c3_7af6;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2795_c3_4584 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2795_c3_4584;
     VAR_sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_y := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2820_c3_47e7 := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2820_c3_47e7;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_72b9_right := to_unsigned(5, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2819_c11_f6eb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_72b9_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue := VAR_previous_stack_read;
     VAR_t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse := t16_high;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse := t16_low;
     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2790_c2_d3ad] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2790_c2_d3ad_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2803_l2806_DUPLICATE_f768 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2803_l2806_DUPLICATE_f768_return_output := result.is_stack_write;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2823_c7_c9e1] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2823_c7_c9e1_return_output := result.stack_address_sp_offset;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2790_c2_d3ad] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2790_c2_d3ad_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l2813_c11_8072] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072_left;
     BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072_return_output := BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2803_l2823_l2790_DUPLICATE_c360 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2803_l2823_l2790_DUPLICATE_c360_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2819_c11_f6eb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2819_c11_f6eb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2819_c11_f6eb_left;
     BIN_OP_EQ_uxn_opcodes_h_l2819_c11_f6eb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2819_c11_f6eb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2819_c11_f6eb_return_output := BIN_OP_EQ_uxn_opcodes_h_l2819_c11_f6eb_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2823_c11_72b9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2823_c11_72b9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_72b9_left;
     BIN_OP_EQ_uxn_opcodes_h_l2823_c11_72b9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_72b9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_72b9_return_output := BIN_OP_EQ_uxn_opcodes_h_l2823_c11_72b9_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2803_l2813_DUPLICATE_db7f LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2803_l2813_DUPLICATE_db7f_return_output := result.sp_relative_shift;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2790_c2_d3ad] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2790_c2_d3ad_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2819_l2813_l2806_l2803_l2823_DUPLICATE_1f5c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2819_l2813_l2806_l2803_l2823_DUPLICATE_1f5c_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2790_c6_3167] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_left;
     BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_return_output := BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2806_c11_aefa] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_left;
     BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_return_output := BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2790_c2_d3ad] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2790_c2_d3ad_return_output := result.is_stack_index_flipped;

     -- sp_relative_shift[uxn_opcodes_h_l2808_c30_ca18] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_ins;
     sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_x;
     sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_return_output := sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2803_c11_0552] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_left;
     BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_return_output := BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_3167_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_0552_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_aefa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_8072_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2819_c11_f6eb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2819_c11_f6eb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2819_c11_f6eb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_72b9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_72b9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_72b9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2803_l2813_DUPLICATE_db7f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2803_l2813_DUPLICATE_db7f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2819_l2813_l2806_l2803_l2823_DUPLICATE_1f5c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2819_l2813_l2806_l2803_l2823_DUPLICATE_1f5c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2819_l2813_l2806_l2803_l2823_DUPLICATE_1f5c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2819_l2813_l2806_l2803_l2823_DUPLICATE_1f5c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2819_l2813_l2806_l2803_l2823_DUPLICATE_1f5c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2803_l2806_DUPLICATE_f768_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2803_l2806_DUPLICATE_f768_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2803_l2823_l2790_DUPLICATE_c360_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2803_l2823_l2790_DUPLICATE_c360_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2803_l2823_l2790_DUPLICATE_c360_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2790_c2_d3ad_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2790_c2_d3ad_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2790_c2_d3ad_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2790_c2_d3ad_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2823_c7_c9e1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2808_c30_ca18_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2813_c7_63d9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2790_c2_d3ad] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2823_c7_c9e1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2790_c2_d3ad] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2790_c2_d3ad] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2823_c7_c9e1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_return_output := result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2790_c2_d3ad] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2806_c7_c4ed] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2806_c7_c4ed] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond;
     t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output := t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2813_c7_63d9] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_cond;
     t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output := t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2823_c7_c9e1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_c9e1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_c9e1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_c9e1_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output;
     -- t16_high_MUX[uxn_opcodes_h_l2803_c7_97e8] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_cond;
     t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output := t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2806_c7_c4ed] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2819_c7_5956] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2819_c7_5956] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_return_output := result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2819_c7_5956] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2806_c7_c4ed] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond;
     t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output := t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2803_c7_97e8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_5956_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_5956_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2819_c7_5956_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2803_c7_97e8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2803_c7_97e8] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_cond;
     t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output := t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2813_c7_63d9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output := result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2813_c7_63d9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2813_c7_63d9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2790_c2_d3ad] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2790_c2_d3ad] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond;
     t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output := t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2813_c7_63d9_return_output;
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2806_c7_c4ed] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2806_c7_c4ed] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2790_c2_d3ad] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2806_c7_c4ed] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output := result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2790_c2_d3ad] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond;
     t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output := t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2806_c7_c4ed_return_output;
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2803_c7_97e8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output := result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2803_c7_97e8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2803_c7_97e8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2803_c7_97e8_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2790_c2_d3ad] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2790_c2_d3ad] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2790_c2_d3ad] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output := result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2829_l2786_DUPLICATE_f68a LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2829_l2786_DUPLICATE_f68a_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8b52(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2790_c2_d3ad_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2829_l2786_DUPLICATE_f68a_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2829_l2786_DUPLICATE_f68a_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
