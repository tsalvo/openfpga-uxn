-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity equ_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end equ_0CLK_226c8821;
architecture arch of equ_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1180_c6_30b6]
signal BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1180_c2_2e6f]
signal t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1180_c2_2e6f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1180_c2_2e6f]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1180_c2_2e6f]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1180_c2_2e6f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1180_c2_2e6f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1180_c2_2e6f]
signal result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1180_c2_2e6f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1180_c2_2e6f]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1180_c2_2e6f]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1180_c2_2e6f]
signal n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1193_c11_344f]
signal BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1193_c7_a491]
signal t8_MUX_uxn_opcodes_h_l1193_c7_a491_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1193_c7_a491_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1193_c7_a491]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1193_c7_a491]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1193_c7_a491]
signal result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1193_c7_a491]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1193_c7_a491]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l1193_c7_a491]
signal n8_MUX_uxn_opcodes_h_l1193_c7_a491_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1193_c7_a491_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1196_c11_e877]
signal BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1196_c7_2fda]
signal t8_MUX_uxn_opcodes_h_l1196_c7_2fda_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1196_c7_2fda]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1196_c7_2fda]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1196_c7_2fda]
signal result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1196_c7_2fda]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1196_c7_2fda]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l1196_c7_2fda]
signal n8_MUX_uxn_opcodes_h_l1196_c7_2fda_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1199_c11_dc8e]
signal BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1199_c7_dfac]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1199_c7_dfac]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1199_c7_dfac]
signal result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1199_c7_dfac]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1199_c7_dfac]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l1199_c7_dfac]
signal n8_MUX_uxn_opcodes_h_l1199_c7_dfac_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1201_c30_12b6]
signal sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1204_c21_3742]
signal BIN_OP_EQ_uxn_opcodes_h_l1204_c21_3742_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1204_c21_3742_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1204_c21_3742_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1204_c21_1d08]
signal MUX_uxn_opcodes_h_l1204_c21_1d08_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1204_c21_1d08_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1204_c21_1d08_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1204_c21_1d08_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c580( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.u8_value := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_stack_index_flipped := ref_toks_8;
      base.is_pc_updated := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6
BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_left,
BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_right,
BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_return_output);

-- t8_MUX_uxn_opcodes_h_l1180_c2_2e6f
t8_MUX_uxn_opcodes_h_l1180_c2_2e6f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond,
t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue,
t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse,
t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f
result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f
result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f
result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f
result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f
result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f
result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output);

-- n8_MUX_uxn_opcodes_h_l1180_c2_2e6f
n8_MUX_uxn_opcodes_h_l1180_c2_2e6f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond,
n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue,
n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse,
n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f
BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_left,
BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_right,
BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_return_output);

-- t8_MUX_uxn_opcodes_h_l1193_c7_a491
t8_MUX_uxn_opcodes_h_l1193_c7_a491 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1193_c7_a491_cond,
t8_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue,
t8_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse,
t8_MUX_uxn_opcodes_h_l1193_c7_a491_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491
result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491
result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_cond,
result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491
result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491
result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_return_output);

-- n8_MUX_uxn_opcodes_h_l1193_c7_a491
n8_MUX_uxn_opcodes_h_l1193_c7_a491 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1193_c7_a491_cond,
n8_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue,
n8_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse,
n8_MUX_uxn_opcodes_h_l1193_c7_a491_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877
BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_left,
BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_right,
BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_return_output);

-- t8_MUX_uxn_opcodes_h_l1196_c7_2fda
t8_MUX_uxn_opcodes_h_l1196_c7_2fda : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1196_c7_2fda_cond,
t8_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue,
t8_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse,
t8_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda
result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda
result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_cond,
result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda
result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda
result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output);

-- n8_MUX_uxn_opcodes_h_l1196_c7_2fda
n8_MUX_uxn_opcodes_h_l1196_c7_2fda : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1196_c7_2fda_cond,
n8_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue,
n8_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse,
n8_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e
BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e_left,
BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e_right,
BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac
result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_cond,
result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac
result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output);

-- n8_MUX_uxn_opcodes_h_l1199_c7_dfac
n8_MUX_uxn_opcodes_h_l1199_c7_dfac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1199_c7_dfac_cond,
n8_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue,
n8_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse,
n8_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6
sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_ins,
sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_x,
sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_y,
sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1204_c21_3742
BIN_OP_EQ_uxn_opcodes_h_l1204_c21_3742 : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1204_c21_3742_left,
BIN_OP_EQ_uxn_opcodes_h_l1204_c21_3742_right,
BIN_OP_EQ_uxn_opcodes_h_l1204_c21_3742_return_output);

-- MUX_uxn_opcodes_h_l1204_c21_1d08
MUX_uxn_opcodes_h_l1204_c21_1d08 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1204_c21_1d08_cond,
MUX_uxn_opcodes_h_l1204_c21_1d08_iftrue,
MUX_uxn_opcodes_h_l1204_c21_1d08_iffalse,
MUX_uxn_opcodes_h_l1204_c21_1d08_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_return_output,
 t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output,
 n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_return_output,
 t8_MUX_uxn_opcodes_h_l1193_c7_a491_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_return_output,
 n8_MUX_uxn_opcodes_h_l1193_c7_a491_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_return_output,
 t8_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output,
 n8_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output,
 n8_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output,
 sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1204_c21_3742_return_output,
 MUX_uxn_opcodes_h_l1204_c21_1d08_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1193_c7_a491_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1180_c2_2e6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1180_c2_2e6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1190_c3_b59a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1185_c3_71c1 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1180_c2_2e6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1180_c2_2e6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1193_c7_a491_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1193_c7_a491_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1194_c3_c417 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1193_c7_a491_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1196_c7_2fda_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1196_c7_2fda_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1203_c3_f86c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1199_c7_dfac_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1204_c21_1d08_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1204_c21_3742_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1204_c21_3742_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1204_c21_3742_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1204_c21_1d08_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1204_c21_1d08_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1204_c21_1d08_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1196_l1180_l1199_l1193_DUPLICATE_6ce3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1196_l1199_l1193_DUPLICATE_3d17_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1196_l1199_l1193_DUPLICATE_7579_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1196_l1199_l1193_DUPLICATE_7c54_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1196_l1199_DUPLICATE_932b_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l1208_l1176_DUPLICATE_8909_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1190_c3_b59a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1190_c3_b59a;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1194_c3_c417 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1194_c3_c417;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1185_c3_71c1 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1185_c3_71c1;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1203_c3_f86c := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1203_c3_f86c;
     VAR_MUX_uxn_opcodes_h_l1204_c21_1d08_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_MUX_uxn_opcodes_h_l1204_c21_1d08_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1204_c21_3742_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1204_c21_3742_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1196_l1199_l1193_DUPLICATE_7579 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1196_l1199_l1193_DUPLICATE_7579_return_output := result.is_stack_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1196_l1199_l1193_DUPLICATE_7c54 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1196_l1199_l1193_DUPLICATE_7c54_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1204_c21_3742] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1204_c21_3742_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1204_c21_3742_left;
     BIN_OP_EQ_uxn_opcodes_h_l1204_c21_3742_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1204_c21_3742_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1204_c21_3742_return_output := BIN_OP_EQ_uxn_opcodes_h_l1204_c21_3742_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1180_c2_2e6f] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1180_c2_2e6f_return_output := result.is_vram_write;

     -- sp_relative_shift[uxn_opcodes_h_l1201_c30_12b6] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_ins;
     sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_x;
     sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_return_output := sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1196_l1199_DUPLICATE_932b LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1196_l1199_DUPLICATE_932b_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1180_c6_30b6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_left;
     BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_return_output := BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1199_c11_dc8e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1193_c11_344f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1180_c2_2e6f] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1180_c2_2e6f_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1196_l1199_l1193_DUPLICATE_3d17 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1196_l1199_l1193_DUPLICATE_3d17_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1196_l1180_l1199_l1193_DUPLICATE_6ce3 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1196_l1180_l1199_l1193_DUPLICATE_6ce3_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1196_c11_e877] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_left;
     BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_return_output := BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1180_c2_2e6f] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1180_c2_2e6f_return_output := result.is_ram_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1180_c2_2e6f] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1180_c2_2e6f_return_output := result.is_pc_updated;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1180_c6_30b6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1193_c7_a491_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1193_c7_a491_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_344f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1196_c7_2fda_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1196_c7_2fda_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_e877_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1199_c7_dfac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_dc8e_return_output;
     VAR_MUX_uxn_opcodes_h_l1204_c21_1d08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1204_c21_3742_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1196_l1199_l1193_DUPLICATE_7c54_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1196_l1199_l1193_DUPLICATE_7c54_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1196_l1199_l1193_DUPLICATE_7c54_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1196_l1199_l1193_DUPLICATE_3d17_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1196_l1199_l1193_DUPLICATE_3d17_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1196_l1199_l1193_DUPLICATE_3d17_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1196_l1199_l1193_DUPLICATE_7579_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1196_l1199_l1193_DUPLICATE_7579_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1196_l1199_l1193_DUPLICATE_7579_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1196_l1199_DUPLICATE_932b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1196_l1199_DUPLICATE_932b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1196_l1180_l1199_l1193_DUPLICATE_6ce3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1196_l1180_l1199_l1193_DUPLICATE_6ce3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1196_l1180_l1199_l1193_DUPLICATE_6ce3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1196_l1180_l1199_l1193_DUPLICATE_6ce3_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1180_c2_2e6f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1180_c2_2e6f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1180_c2_2e6f_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1180_c2_2e6f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1201_c30_12b6_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1199_c7_dfac] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output;

     -- MUX[uxn_opcodes_h_l1204_c21_1d08] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1204_c21_1d08_cond <= VAR_MUX_uxn_opcodes_h_l1204_c21_1d08_cond;
     MUX_uxn_opcodes_h_l1204_c21_1d08_iftrue <= VAR_MUX_uxn_opcodes_h_l1204_c21_1d08_iftrue;
     MUX_uxn_opcodes_h_l1204_c21_1d08_iffalse <= VAR_MUX_uxn_opcodes_h_l1204_c21_1d08_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1204_c21_1d08_return_output := MUX_uxn_opcodes_h_l1204_c21_1d08_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1180_c2_2e6f] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output;

     -- t8_MUX[uxn_opcodes_h_l1196_c7_2fda] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1196_c7_2fda_cond <= VAR_t8_MUX_uxn_opcodes_h_l1196_c7_2fda_cond;
     t8_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue;
     t8_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output := t8_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1199_c7_dfac] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output;

     -- n8_MUX[uxn_opcodes_h_l1199_c7_dfac] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1199_c7_dfac_cond <= VAR_n8_MUX_uxn_opcodes_h_l1199_c7_dfac_cond;
     n8_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue;
     n8_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output := n8_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1180_c2_2e6f] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1180_c2_2e6f] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1199_c7_dfac] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1199_c7_dfac] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1180_c2_2e6f] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue := VAR_MUX_uxn_opcodes_h_l1204_c21_1d08_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1196_c7_2fda] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1196_c7_2fda] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output;

     -- t8_MUX[uxn_opcodes_h_l1193_c7_a491] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1193_c7_a491_cond <= VAR_t8_MUX_uxn_opcodes_h_l1193_c7_a491_cond;
     t8_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue;
     t8_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1193_c7_a491_return_output := t8_MUX_uxn_opcodes_h_l1193_c7_a491_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1199_c7_dfac] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output := result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1196_c7_2fda] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1196_c7_2fda] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output;

     -- n8_MUX[uxn_opcodes_h_l1196_c7_2fda] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1196_c7_2fda_cond <= VAR_n8_MUX_uxn_opcodes_h_l1196_c7_2fda_cond;
     n8_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue;
     n8_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output := n8_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_dfac_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1193_c7_a491_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1193_c7_a491] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1193_c7_a491] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_return_output;

     -- t8_MUX[uxn_opcodes_h_l1180_c2_2e6f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond <= VAR_t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond;
     t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue;
     t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output := t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output;

     -- n8_MUX[uxn_opcodes_h_l1193_c7_a491] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1193_c7_a491_cond <= VAR_n8_MUX_uxn_opcodes_h_l1193_c7_a491_cond;
     n8_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue;
     n8_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1193_c7_a491_return_output := n8_MUX_uxn_opcodes_h_l1193_c7_a491_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1193_c7_a491] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1193_c7_a491] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1196_c7_2fda] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output := result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1193_c7_a491_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_a491_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_a491_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_a491_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_a491_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_2fda_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1193_c7_a491] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_return_output := result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1180_c2_2e6f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1180_c2_2e6f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1180_c2_2e6f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output;

     -- n8_MUX[uxn_opcodes_h_l1180_c2_2e6f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond <= VAR_n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond;
     n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue;
     n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output := n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1180_c2_2e6f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_a491_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1180_c2_2e6f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l1208_l1176_DUPLICATE_8909 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l1208_l1176_DUPLICATE_8909_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c580(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1180_c2_2e6f_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l1208_l1176_DUPLICATE_8909_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l1208_l1176_DUPLICATE_8909_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
