-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 56
entity jsr_0CLK_6da26caa is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jsr_0CLK_6da26caa;
architecture arch of jsr_0CLK_6da26caa is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l706_c6_8b1e]
signal BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l706_c1_4926]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l706_c2_d762]
signal t8_MUX_uxn_opcodes_h_l706_c2_d762_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l706_c2_d762_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l706_c2_d762_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l706_c2_d762_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l706_c2_d762]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l706_c2_d762]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l706_c2_d762]
signal result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l706_c2_d762]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l706_c2_d762]
signal result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l706_c2_d762]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l706_c2_d762]
signal result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l706_c2_d762]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l706_c2_d762]
signal result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_return_output : unsigned(15 downto 0);

-- printf_uxn_opcodes_h_l707_c3_70b6[uxn_opcodes_h_l707_c3_70b6]
signal printf_uxn_opcodes_h_l707_c3_70b6_uxn_opcodes_h_l707_c3_70b6_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l711_c11_58b5]
signal BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l711_c7_94b2]
signal t8_MUX_uxn_opcodes_h_l711_c7_94b2_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l711_c7_94b2_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l711_c7_94b2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l711_c7_94b2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l711_c7_94b2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l711_c7_94b2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l711_c7_94b2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l711_c7_94b2]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l711_c7_94b2]
signal result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l711_c7_94b2]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l711_c7_94b2]
signal result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l714_c30_d295]
signal sp_relative_shift_uxn_opcodes_h_l714_c30_d295_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l714_c30_d295_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l714_c30_d295_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l714_c30_d295_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l716_c11_2388]
signal BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l716_c7_bfc4]
signal t8_MUX_uxn_opcodes_h_l716_c7_bfc4_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l716_c7_bfc4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l716_c7_bfc4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l716_c7_bfc4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l716_c7_bfc4]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l716_c7_bfc4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l716_c7_bfc4]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l716_c7_bfc4]
signal result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l716_c7_bfc4]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l716_c7_bfc4]
signal result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l724_c11_503c]
signal BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l724_c7_fd44]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l724_c7_fd44]
signal result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l724_c7_fd44]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l724_c7_fd44]
signal result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l724_c7_fd44]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l724_c7_fd44]
signal result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l724_c7_fd44]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l724_c7_fd44]
signal result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_return_output : unsigned(15 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l727_c31_1266]
signal CONST_SR_8_uxn_opcodes_h_l727_c31_1266_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l727_c31_1266_return_output : unsigned(15 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l729_c22_0fcc]
signal BIN_OP_PLUS_uxn_opcodes_h_l729_c22_0fcc_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l729_c22_0fcc_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l729_c22_0fcc_return_output : signed(17 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l731_c11_1bdd]
signal BIN_OP_EQ_uxn_opcodes_h_l731_c11_1bdd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l731_c11_1bdd_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l731_c11_1bdd_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l731_c7_38c8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l731_c7_38c8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l731_c7_38c8]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l731_c7_38c8]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_return_output : unsigned(0 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_3dbc( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : signed;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.sp_relative_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_sp_shift := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.u16_value := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e
BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_left,
BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_right,
BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_return_output);

-- t8_MUX_uxn_opcodes_h_l706_c2_d762
t8_MUX_uxn_opcodes_h_l706_c2_d762 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l706_c2_d762_cond,
t8_MUX_uxn_opcodes_h_l706_c2_d762_iftrue,
t8_MUX_uxn_opcodes_h_l706_c2_d762_iffalse,
t8_MUX_uxn_opcodes_h_l706_c2_d762_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762
result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762
result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762
result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762
result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762
result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_cond,
result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762
result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762
result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_cond,
result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_return_output);

-- printf_uxn_opcodes_h_l707_c3_70b6_uxn_opcodes_h_l707_c3_70b6
printf_uxn_opcodes_h_l707_c3_70b6_uxn_opcodes_h_l707_c3_70b6 : entity work.printf_uxn_opcodes_h_l707_c3_70b6_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l707_c3_70b6_uxn_opcodes_h_l707_c3_70b6_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5
BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_left,
BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_right,
BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_return_output);

-- t8_MUX_uxn_opcodes_h_l711_c7_94b2
t8_MUX_uxn_opcodes_h_l711_c7_94b2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l711_c7_94b2_cond,
t8_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue,
t8_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse,
t8_MUX_uxn_opcodes_h_l711_c7_94b2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2
result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2
result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2
result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2
result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2
result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_cond,
result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2
result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2
result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_cond,
result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_return_output);

-- sp_relative_shift_uxn_opcodes_h_l714_c30_d295
sp_relative_shift_uxn_opcodes_h_l714_c30_d295 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l714_c30_d295_ins,
sp_relative_shift_uxn_opcodes_h_l714_c30_d295_x,
sp_relative_shift_uxn_opcodes_h_l714_c30_d295_y,
sp_relative_shift_uxn_opcodes_h_l714_c30_d295_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388
BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_left,
BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_right,
BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_return_output);

-- t8_MUX_uxn_opcodes_h_l716_c7_bfc4
t8_MUX_uxn_opcodes_h_l716_c7_bfc4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l716_c7_bfc4_cond,
t8_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue,
t8_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse,
t8_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4
result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4
result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4
result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4
result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4
result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_cond,
result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4
result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4
result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_cond,
result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c
BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_left,
BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_right,
BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44
result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44
result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44
result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44
result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_cond,
result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44
result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44
result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_cond,
result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_return_output);

-- CONST_SR_8_uxn_opcodes_h_l727_c31_1266
CONST_SR_8_uxn_opcodes_h_l727_c31_1266 : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l727_c31_1266_x,
CONST_SR_8_uxn_opcodes_h_l727_c31_1266_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l729_c22_0fcc
BIN_OP_PLUS_uxn_opcodes_h_l729_c22_0fcc : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l729_c22_0fcc_left,
BIN_OP_PLUS_uxn_opcodes_h_l729_c22_0fcc_right,
BIN_OP_PLUS_uxn_opcodes_h_l729_c22_0fcc_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l731_c11_1bdd
BIN_OP_EQ_uxn_opcodes_h_l731_c11_1bdd : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l731_c11_1bdd_left,
BIN_OP_EQ_uxn_opcodes_h_l731_c11_1bdd_right,
BIN_OP_EQ_uxn_opcodes_h_l731_c11_1bdd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8
result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8
result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8
result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_return_output,
 t8_MUX_uxn_opcodes_h_l706_c2_d762_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_return_output,
 t8_MUX_uxn_opcodes_h_l711_c7_94b2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_return_output,
 sp_relative_shift_uxn_opcodes_h_l714_c30_d295_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_return_output,
 t8_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_return_output,
 CONST_SR_8_uxn_opcodes_h_l727_c31_1266_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l729_c22_0fcc_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l731_c11_1bdd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l706_c2_d762_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l706_c2_d762_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l711_c7_94b2_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l706_c2_d762_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l706_c2_d762_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l708_c3_c46a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l707_c3_70b6_uxn_opcodes_h_l707_c3_70b6_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l711_c7_94b2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l712_c3_aa34 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l714_c30_d295_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l714_c30_d295_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l714_c30_d295_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l714_c30_d295_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l716_c7_bfc4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l721_c3_7373 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l719_c3_3f4e : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_cond : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l722_c21_59ad_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l726_c3_3bbe : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l724_c7_fd44_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l729_c3_b342 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l727_c31_1266_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l727_c31_1266_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l727_c21_ee69_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l729_c22_0fcc_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l729_c27_59a7_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l729_c22_0fcc_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l729_c22_0fcc_return_output : signed(17 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l731_c11_1bdd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l731_c11_1bdd_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l731_c11_1bdd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l716_l706_DUPLICATE_c50f_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l716_l706_l724_DUPLICATE_3e5d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l711_l731_l706_l724_DUPLICATE_59cc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l711_l731_l706_l724_DUPLICATE_fd53_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l711_l706_l724_DUPLICATE_f25b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l711_l731_l716_l706_DUPLICATE_6f91_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l711_l716_l706_l724_DUPLICATE_93ab_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l711_l731_l716_l724_DUPLICATE_ef66_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3dbc_uxn_opcodes_h_l738_l702_DUPLICATE_02e3_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l726_c3_3bbe := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l726_c3_3bbe;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l712_c3_aa34 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l712_c3_aa34;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l714_c30_d295_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_right := to_unsigned(3, 2);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_iffalse := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l714_c30_d295_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l708_c3_c46a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l708_c3_c46a;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l731_c11_1bdd_right := to_unsigned(4, 3);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l719_c3_3f4e := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l719_c3_3f4e;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l721_c3_7373 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l721_c3_7373;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l714_c30_d295_ins := VAR_ins;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l729_c22_0fcc_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_CONST_SR_8_uxn_opcodes_h_l727_c31_1266_x := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l731_c11_1bdd_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l706_c2_d762_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l711_l731_l716_l724_DUPLICATE_ef66 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l711_l731_l716_l724_DUPLICATE_ef66_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l711_c11_58b5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_left;
     BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_return_output := BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l711_l731_l706_l724_DUPLICATE_59cc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l711_l731_l706_l724_DUPLICATE_59cc_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l711_l731_l706_l724_DUPLICATE_fd53 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l711_l731_l706_l724_DUPLICATE_fd53_return_output := result.is_stack_index_flipped;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l722_c21_59ad] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l722_c21_59ad_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_pc);

     -- CAST_TO_int8_t[uxn_opcodes_h_l729_c27_59a7] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l729_c27_59a7_return_output := CAST_TO_int8_t_uint8_t(
     t8);

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l711_l716_l706_l724_DUPLICATE_93ab LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l711_l716_l706_l724_DUPLICATE_93ab_return_output := result.u16_value;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l724_c7_fd44] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l724_c7_fd44_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l706_c6_8b1e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_left;
     BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_return_output := BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l724_c11_503c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_left;
     BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_return_output := BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_return_output;

     -- CONST_SR_8[uxn_opcodes_h_l727_c31_1266] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l727_c31_1266_x <= VAR_CONST_SR_8_uxn_opcodes_h_l727_c31_1266_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l727_c31_1266_return_output := CONST_SR_8_uxn_opcodes_h_l727_c31_1266_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l731_c11_1bdd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l731_c11_1bdd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l731_c11_1bdd_left;
     BIN_OP_EQ_uxn_opcodes_h_l731_c11_1bdd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l731_c11_1bdd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l731_c11_1bdd_return_output := BIN_OP_EQ_uxn_opcodes_h_l731_c11_1bdd_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l711_l731_l716_l706_DUPLICATE_6f91 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l711_l731_l716_l706_DUPLICATE_6f91_return_output := result.is_pc_updated;

     -- sp_relative_shift[uxn_opcodes_h_l714_c30_d295] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l714_c30_d295_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l714_c30_d295_ins;
     sp_relative_shift_uxn_opcodes_h_l714_c30_d295_x <= VAR_sp_relative_shift_uxn_opcodes_h_l714_c30_d295_x;
     sp_relative_shift_uxn_opcodes_h_l714_c30_d295_y <= VAR_sp_relative_shift_uxn_opcodes_h_l714_c30_d295_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l714_c30_d295_return_output := sp_relative_shift_uxn_opcodes_h_l714_c30_d295_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l716_c11_2388] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_left;
     BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_return_output := BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l716_l706_DUPLICATE_c50f LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l716_l706_DUPLICATE_c50f_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l716_l706_l724_DUPLICATE_3e5d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l716_l706_l724_DUPLICATE_3e5d_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l711_l706_l724_DUPLICATE_f25b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l711_l706_l724_DUPLICATE_f25b_return_output := result.u8_value;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l706_c2_d762_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c6_8b1e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l711_c7_94b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l711_c11_58b5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l716_c7_bfc4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l716_c11_2388_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l724_c11_503c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l731_c11_1bdd_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l731_c11_1bdd_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l731_c11_1bdd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l731_c11_1bdd_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l729_c22_0fcc_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l729_c27_59a7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l722_c21_59ad_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l716_l706_DUPLICATE_c50f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l716_l706_DUPLICATE_c50f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l711_l716_l706_l724_DUPLICATE_93ab_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l711_l716_l706_l724_DUPLICATE_93ab_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l711_l716_l706_l724_DUPLICATE_93ab_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l711_l716_l706_l724_DUPLICATE_93ab_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l711_l731_l716_l724_DUPLICATE_ef66_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l711_l731_l716_l724_DUPLICATE_ef66_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l711_l731_l716_l724_DUPLICATE_ef66_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l711_l731_l716_l724_DUPLICATE_ef66_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l711_l731_l716_l706_DUPLICATE_6f91_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l711_l731_l716_l706_DUPLICATE_6f91_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l711_l731_l716_l706_DUPLICATE_6f91_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l711_l731_l716_l706_DUPLICATE_6f91_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l716_l706_l724_DUPLICATE_3e5d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l716_l706_l724_DUPLICATE_3e5d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l716_l706_l724_DUPLICATE_3e5d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l711_l731_l706_l724_DUPLICATE_fd53_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l711_l731_l706_l724_DUPLICATE_fd53_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l711_l731_l706_l724_DUPLICATE_fd53_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l711_l731_l706_l724_DUPLICATE_fd53_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l711_l731_l706_l724_DUPLICATE_59cc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l711_l731_l706_l724_DUPLICATE_59cc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l711_l731_l706_l724_DUPLICATE_59cc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l711_l731_l706_l724_DUPLICATE_59cc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l711_l706_l724_DUPLICATE_f25b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l711_l706_l724_DUPLICATE_f25b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l711_l706_l724_DUPLICATE_f25b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l724_c7_fd44_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l714_c30_d295_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l706_c1_4926] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l727_c21_ee69] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l727_c21_ee69_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l727_c31_1266_return_output);

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l724_c7_fd44] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l724_c7_fd44] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l731_c7_38c8] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l731_c7_38c8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l716_c7_bfc4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l731_c7_38c8] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l729_c22_0fcc] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l729_c22_0fcc_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l729_c22_0fcc_left;
     BIN_OP_PLUS_uxn_opcodes_h_l729_c22_0fcc_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l729_c22_0fcc_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l729_c22_0fcc_return_output := BIN_OP_PLUS_uxn_opcodes_h_l729_c22_0fcc_return_output;

     -- t8_MUX[uxn_opcodes_h_l716_c7_bfc4] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l716_c7_bfc4_cond <= VAR_t8_MUX_uxn_opcodes_h_l716_c7_bfc4_cond;
     t8_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue;
     t8_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output := t8_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l731_c7_38c8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_return_output;

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l729_c3_b342 := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l729_c22_0fcc_return_output)),16);
     VAR_result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l727_c21_ee69_return_output;
     VAR_printf_uxn_opcodes_h_l707_c3_70b6_uxn_opcodes_h_l707_c3_70b6_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l706_c1_4926_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l731_c7_38c8_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l731_c7_38c8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l724_c7_fd44_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l731_c7_38c8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l731_c7_38c8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l724_c7_fd44_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse := VAR_t8_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue := VAR_result_u16_value_uxn_opcodes_h_l729_c3_b342;
     -- t8_MUX[uxn_opcodes_h_l711_c7_94b2] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l711_c7_94b2_cond <= VAR_t8_MUX_uxn_opcodes_h_l711_c7_94b2_cond;
     t8_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue;
     t8_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l711_c7_94b2_return_output := t8_MUX_uxn_opcodes_h_l711_c7_94b2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l716_c7_bfc4] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l724_c7_fd44] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l724_c7_fd44] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_cond;
     result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_return_output := result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l716_c7_bfc4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l724_c7_fd44] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l724_c7_fd44] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l711_c7_94b2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l724_c7_fd44] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_return_output;

     -- printf_uxn_opcodes_h_l707_c3_70b6[uxn_opcodes_h_l707_c3_70b6] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l707_c3_70b6_uxn_opcodes_h_l707_c3_70b6_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l707_c3_70b6_uxn_opcodes_h_l707_c3_70b6_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_u8_value_MUX[uxn_opcodes_h_l724_c7_fd44] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_cond;
     result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_return_output := result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l724_c7_fd44_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l724_c7_fd44_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l724_c7_fd44_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l724_c7_fd44_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l711_c7_94b2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l724_c7_fd44_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l724_c7_fd44_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l706_c2_d762_iffalse := VAR_t8_MUX_uxn_opcodes_h_l711_c7_94b2_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l716_c7_bfc4] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_cond;
     result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output := result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l706_c2_d762] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l711_c7_94b2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l716_c7_bfc4] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l716_c7_bfc4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output;

     -- t8_MUX[uxn_opcodes_h_l706_c2_d762] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l706_c2_d762_cond <= VAR_t8_MUX_uxn_opcodes_h_l706_c2_d762_cond;
     t8_MUX_uxn_opcodes_h_l706_c2_d762_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l706_c2_d762_iftrue;
     t8_MUX_uxn_opcodes_h_l706_c2_d762_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l706_c2_d762_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l706_c2_d762_return_output := t8_MUX_uxn_opcodes_h_l706_c2_d762_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l716_c7_bfc4] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l716_c7_bfc4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l711_c7_94b2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l716_c7_bfc4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output := result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l711_c7_94b2_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l711_c7_94b2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l716_c7_bfc4_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l706_c2_d762_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l711_c7_94b2] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l711_c7_94b2] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l711_c7_94b2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l706_c2_d762] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l711_c7_94b2] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_cond;
     result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_return_output := result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l711_c7_94b2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_return_output := result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l706_c2_d762] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l711_c7_94b2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l711_c7_94b2_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l711_c7_94b2_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l711_c7_94b2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l711_c7_94b2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l711_c7_94b2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l711_c7_94b2_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l706_c2_d762] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l706_c2_d762] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_cond;
     result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_return_output := result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l706_c2_d762] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l706_c2_d762] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_cond;
     result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_return_output := result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l706_c2_d762] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l706_c2_d762] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_3dbc_uxn_opcodes_h_l738_l702_DUPLICATE_02e3 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3dbc_uxn_opcodes_h_l738_l702_DUPLICATE_02e3_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_3dbc(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l706_c2_d762_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l706_c2_d762_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l706_c2_d762_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l706_c2_d762_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l706_c2_d762_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l706_c2_d762_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l706_c2_d762_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l706_c2_d762_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l706_c2_d762_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3dbc_uxn_opcodes_h_l738_l702_DUPLICATE_02e3_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3dbc_uxn_opcodes_h_l738_l702_DUPLICATE_02e3_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
