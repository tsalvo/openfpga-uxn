-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 52
entity ora_0CLK_f62d646e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ora_0CLK_f62d646e;
architecture arch of ora_0CLK_f62d646e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1045_c6_b1d2]
signal BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1045_c1_e619]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1045_c2_548e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1045_c2_548e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1045_c2_548e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1045_c2_548e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1045_c2_548e]
signal result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1045_c2_548e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1045_c2_548e]
signal t8_MUX_uxn_opcodes_h_l1045_c2_548e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1045_c2_548e_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1045_c2_548e]
signal n8_MUX_uxn_opcodes_h_l1045_c2_548e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1045_c2_548e_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1046_c3_53ee[uxn_opcodes_h_l1046_c3_53ee]
signal printf_uxn_opcodes_h_l1046_c3_53ee_uxn_opcodes_h_l1046_c3_53ee_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1050_c11_bd91]
signal BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1050_c7_eab2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1050_c7_eab2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1050_c7_eab2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1050_c7_eab2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1050_c7_eab2]
signal result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1050_c7_eab2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1050_c7_eab2]
signal t8_MUX_uxn_opcodes_h_l1050_c7_eab2_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1050_c7_eab2]
signal n8_MUX_uxn_opcodes_h_l1050_c7_eab2_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1053_c11_640b]
signal BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1053_c7_4fa5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1053_c7_4fa5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1053_c7_4fa5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1053_c7_4fa5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1053_c7_4fa5]
signal result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1053_c7_4fa5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1053_c7_4fa5]
signal t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1053_c7_4fa5]
signal n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1057_c11_79ca]
signal BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1057_c7_6bed]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1057_c7_6bed]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1057_c7_6bed]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1057_c7_6bed]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1057_c7_6bed]
signal result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1057_c7_6bed]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l1057_c7_6bed]
signal n8_MUX_uxn_opcodes_h_l1057_c7_6bed_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1060_c11_9f66]
signal BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1060_c7_94d2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1060_c7_94d2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1060_c7_94d2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1060_c7_94d2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1060_c7_94d2]
signal result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1060_c7_94d2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l1060_c7_94d2]
signal n8_MUX_uxn_opcodes_h_l1060_c7_94d2_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1063_c30_2624]
signal sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_return_output : signed(3 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l1066_c21_8ecf]
signal BIN_OP_OR_uxn_opcodes_h_l1066_c21_8ecf_left : unsigned(7 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l1066_c21_8ecf_right : unsigned(7 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l1066_c21_8ecf_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1068_c11_60bd]
signal BIN_OP_EQ_uxn_opcodes_h_l1068_c11_60bd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1068_c11_60bd_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1068_c11_60bd_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1068_c7_237f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1068_c7_237f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1068_c7_237f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_641b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2
BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_left,
BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_right,
BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e
result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e
result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e
result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e
result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_cond,
result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e
result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_return_output);

-- t8_MUX_uxn_opcodes_h_l1045_c2_548e
t8_MUX_uxn_opcodes_h_l1045_c2_548e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1045_c2_548e_cond,
t8_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue,
t8_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse,
t8_MUX_uxn_opcodes_h_l1045_c2_548e_return_output);

-- n8_MUX_uxn_opcodes_h_l1045_c2_548e
n8_MUX_uxn_opcodes_h_l1045_c2_548e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1045_c2_548e_cond,
n8_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue,
n8_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse,
n8_MUX_uxn_opcodes_h_l1045_c2_548e_return_output);

-- printf_uxn_opcodes_h_l1046_c3_53ee_uxn_opcodes_h_l1046_c3_53ee
printf_uxn_opcodes_h_l1046_c3_53ee_uxn_opcodes_h_l1046_c3_53ee : entity work.printf_uxn_opcodes_h_l1046_c3_53ee_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1046_c3_53ee_uxn_opcodes_h_l1046_c3_53ee_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91
BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_left,
BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_right,
BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2
result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2
result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2
result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2
result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_cond,
result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2
result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output);

-- t8_MUX_uxn_opcodes_h_l1050_c7_eab2
t8_MUX_uxn_opcodes_h_l1050_c7_eab2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1050_c7_eab2_cond,
t8_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue,
t8_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse,
t8_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output);

-- n8_MUX_uxn_opcodes_h_l1050_c7_eab2
n8_MUX_uxn_opcodes_h_l1050_c7_eab2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1050_c7_eab2_cond,
n8_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue,
n8_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse,
n8_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b
BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_left,
BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_right,
BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5
result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5
result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5
result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5
result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond,
result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5
result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output);

-- t8_MUX_uxn_opcodes_h_l1053_c7_4fa5
t8_MUX_uxn_opcodes_h_l1053_c7_4fa5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond,
t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue,
t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse,
t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output);

-- n8_MUX_uxn_opcodes_h_l1053_c7_4fa5
n8_MUX_uxn_opcodes_h_l1053_c7_4fa5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond,
n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue,
n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse,
n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca
BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_left,
BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_right,
BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed
result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed
result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed
result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed
result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_cond,
result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed
result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output);

-- n8_MUX_uxn_opcodes_h_l1057_c7_6bed
n8_MUX_uxn_opcodes_h_l1057_c7_6bed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1057_c7_6bed_cond,
n8_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue,
n8_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse,
n8_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66
BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_left,
BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_right,
BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2
result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2
result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2
result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2
result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_cond,
result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2
result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output);

-- n8_MUX_uxn_opcodes_h_l1060_c7_94d2
n8_MUX_uxn_opcodes_h_l1060_c7_94d2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1060_c7_94d2_cond,
n8_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue,
n8_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse,
n8_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1063_c30_2624
sp_relative_shift_uxn_opcodes_h_l1063_c30_2624 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_ins,
sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_x,
sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_y,
sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l1066_c21_8ecf
BIN_OP_OR_uxn_opcodes_h_l1066_c21_8ecf : entity work.BIN_OP_OR_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l1066_c21_8ecf_left,
BIN_OP_OR_uxn_opcodes_h_l1066_c21_8ecf_right,
BIN_OP_OR_uxn_opcodes_h_l1066_c21_8ecf_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1068_c11_60bd
BIN_OP_EQ_uxn_opcodes_h_l1068_c11_60bd : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1068_c11_60bd_left,
BIN_OP_EQ_uxn_opcodes_h_l1068_c11_60bd_right,
BIN_OP_EQ_uxn_opcodes_h_l1068_c11_60bd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f
result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f
result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f
result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_return_output,
 t8_MUX_uxn_opcodes_h_l1045_c2_548e_return_output,
 n8_MUX_uxn_opcodes_h_l1045_c2_548e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output,
 t8_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output,
 n8_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output,
 t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output,
 n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output,
 n8_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output,
 n8_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output,
 sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_return_output,
 BIN_OP_OR_uxn_opcodes_h_l1066_c21_8ecf_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1068_c11_60bd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_iffalse : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1047_c3_c47b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1045_c2_548e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1045_c2_548e_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1045_c2_548e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1045_c2_548e_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1046_c3_53ee_uxn_opcodes_h_l1046_c3_53ee_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1051_c3_6361 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1050_c7_eab2_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1050_c7_eab2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1055_c3_d0bb : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1058_c3_4a55 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1057_c7_6bed_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1065_c3_cd70 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1060_c7_94d2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1060_c7_94d2_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1066_c21_8ecf_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1066_c21_8ecf_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1066_c21_8ecf_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1068_c11_60bd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1068_c11_60bd_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1068_c11_60bd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1050_l1045_l1068_l1057_l1053_DUPLICATE_8682_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1050_l1045_l1068_l1057_l1053_DUPLICATE_ba41_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1050_l1045_l1060_l1057_l1053_DUPLICATE_a327_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1050_l1045_l1060_l1057_l1053_DUPLICATE_c124_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1050_l1068_l1060_l1057_l1053_DUPLICATE_be93_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1074_l1041_DUPLICATE_34fe_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1068_c11_60bd_right := to_unsigned(5, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1065_c3_cd70 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1065_c3_cd70;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1055_c3_d0bb := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1055_c3_d0bb;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1051_c3_6361 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1051_c3_6361;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1058_c3_4a55 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1058_c3_4a55;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1047_c3_c47b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1047_c3_c47b;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1068_c11_60bd_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l1066_c21_8ecf_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_OR_uxn_opcodes_h_l1066_c21_8ecf_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse := t8;
     -- sp_relative_shift[uxn_opcodes_h_l1063_c30_2624] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_ins;
     sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_x;
     sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_return_output := sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1053_c11_640b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1050_l1045_l1060_l1057_l1053_DUPLICATE_a327 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1050_l1045_l1060_l1057_l1053_DUPLICATE_a327_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1068_c11_60bd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1068_c11_60bd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1068_c11_60bd_left;
     BIN_OP_EQ_uxn_opcodes_h_l1068_c11_60bd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1068_c11_60bd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1068_c11_60bd_return_output := BIN_OP_EQ_uxn_opcodes_h_l1068_c11_60bd_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1050_l1045_l1068_l1057_l1053_DUPLICATE_ba41 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1050_l1045_l1068_l1057_l1053_DUPLICATE_ba41_return_output := result.is_stack_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1050_l1045_l1060_l1057_l1053_DUPLICATE_c124 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1050_l1045_l1060_l1057_l1053_DUPLICATE_c124_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1057_c11_79ca] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_left;
     BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_return_output := BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l1066_c21_8ecf] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l1066_c21_8ecf_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l1066_c21_8ecf_left;
     BIN_OP_OR_uxn_opcodes_h_l1066_c21_8ecf_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l1066_c21_8ecf_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l1066_c21_8ecf_return_output := BIN_OP_OR_uxn_opcodes_h_l1066_c21_8ecf_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1060_c7_94d2] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1060_c7_94d2_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1060_c11_9f66] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_left;
     BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_return_output := BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1050_l1068_l1060_l1057_l1053_DUPLICATE_be93 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1050_l1068_l1060_l1057_l1053_DUPLICATE_be93_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1045_c6_b1d2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_left;
     BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_return_output := BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1050_l1045_l1068_l1057_l1053_DUPLICATE_8682 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1050_l1045_l1068_l1057_l1053_DUPLICATE_8682_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1050_c11_bd91] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_left;
     BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_return_output := BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1045_c2_548e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1045_c2_548e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1045_c6_b1d2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1050_c7_eab2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1050_c7_eab2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1050_c11_bd91_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1053_c11_640b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1057_c7_6bed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1057_c11_79ca_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1060_c7_94d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1060_c11_9f66_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1068_c11_60bd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1068_c11_60bd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1068_c11_60bd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l1066_c21_8ecf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1050_l1045_l1060_l1057_l1053_DUPLICATE_c124_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1050_l1045_l1060_l1057_l1053_DUPLICATE_c124_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1050_l1045_l1060_l1057_l1053_DUPLICATE_c124_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1050_l1045_l1060_l1057_l1053_DUPLICATE_c124_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1050_l1045_l1060_l1057_l1053_DUPLICATE_c124_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1050_l1068_l1060_l1057_l1053_DUPLICATE_be93_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1050_l1068_l1060_l1057_l1053_DUPLICATE_be93_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1050_l1068_l1060_l1057_l1053_DUPLICATE_be93_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1050_l1068_l1060_l1057_l1053_DUPLICATE_be93_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1050_l1068_l1060_l1057_l1053_DUPLICATE_be93_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1050_l1045_l1068_l1057_l1053_DUPLICATE_8682_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1050_l1045_l1068_l1057_l1053_DUPLICATE_8682_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1050_l1045_l1068_l1057_l1053_DUPLICATE_8682_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1050_l1045_l1068_l1057_l1053_DUPLICATE_8682_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1050_l1045_l1068_l1057_l1053_DUPLICATE_8682_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1050_l1045_l1068_l1057_l1053_DUPLICATE_ba41_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1050_l1045_l1068_l1057_l1053_DUPLICATE_ba41_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1050_l1045_l1068_l1057_l1053_DUPLICATE_ba41_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1050_l1045_l1068_l1057_l1053_DUPLICATE_ba41_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1050_l1045_l1068_l1057_l1053_DUPLICATE_ba41_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1050_l1045_l1060_l1057_l1053_DUPLICATE_a327_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1050_l1045_l1060_l1057_l1053_DUPLICATE_a327_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1050_l1045_l1060_l1057_l1053_DUPLICATE_a327_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1050_l1045_l1060_l1057_l1053_DUPLICATE_a327_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1050_l1045_l1060_l1057_l1053_DUPLICATE_a327_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1060_c7_94d2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1063_c30_2624_return_output;
     -- t8_MUX[uxn_opcodes_h_l1053_c7_4fa5] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond <= VAR_t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond;
     t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue;
     t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output := t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1068_c7_237f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1060_c7_94d2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1068_c7_237f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1060_c7_94d2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1068_c7_237f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_return_output;

     -- n8_MUX[uxn_opcodes_h_l1060_c7_94d2] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1060_c7_94d2_cond <= VAR_n8_MUX_uxn_opcodes_h_l1060_c7_94d2_cond;
     n8_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue;
     n8_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output := n8_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1045_c1_e619] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1060_c7_94d2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output := result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l1046_c3_53ee_uxn_opcodes_h_l1046_c3_53ee_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1045_c1_e619_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1068_c7_237f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1068_c7_237f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1068_c7_237f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1057_c7_6bed] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output;

     -- n8_MUX[uxn_opcodes_h_l1057_c7_6bed] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1057_c7_6bed_cond <= VAR_n8_MUX_uxn_opcodes_h_l1057_c7_6bed_cond;
     n8_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue;
     n8_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output := n8_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output;

     -- t8_MUX[uxn_opcodes_h_l1050_c7_eab2] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1050_c7_eab2_cond <= VAR_t8_MUX_uxn_opcodes_h_l1050_c7_eab2_cond;
     t8_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue;
     t8_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output := t8_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1060_c7_94d2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1060_c7_94d2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1057_c7_6bed] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1060_c7_94d2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output;

     -- printf_uxn_opcodes_h_l1046_c3_53ee[uxn_opcodes_h_l1046_c3_53ee] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1046_c3_53ee_uxn_opcodes_h_l1046_c3_53ee_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1046_c3_53ee_uxn_opcodes_h_l1046_c3_53ee_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_u8_value_MUX[uxn_opcodes_h_l1057_c7_6bed] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output := result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1060_c7_94d2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output;
     -- t8_MUX[uxn_opcodes_h_l1045_c2_548e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1045_c2_548e_cond <= VAR_t8_MUX_uxn_opcodes_h_l1045_c2_548e_cond;
     t8_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue;
     t8_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1045_c2_548e_return_output := t8_MUX_uxn_opcodes_h_l1045_c2_548e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1053_c7_4fa5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output := result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1053_c7_4fa5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1057_c7_6bed] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output;

     -- n8_MUX[uxn_opcodes_h_l1053_c7_4fa5] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond <= VAR_n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond;
     n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue;
     n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output := n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1057_c7_6bed] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1053_c7_4fa5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1057_c7_6bed] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1057_c7_6bed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1045_c2_548e_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1050_c7_eab2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1053_c7_4fa5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1050_c7_eab2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output := result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1053_c7_4fa5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1053_c7_4fa5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1050_c7_eab2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output;

     -- n8_MUX[uxn_opcodes_h_l1050_c7_eab2] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1050_c7_eab2_cond <= VAR_n8_MUX_uxn_opcodes_h_l1050_c7_eab2_cond;
     n8_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue;
     n8_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output := n8_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1053_c7_4fa5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1050_c7_eab2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1045_c2_548e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1045_c2_548e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_return_output := result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1050_c7_eab2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1050_c7_eab2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output;

     -- n8_MUX[uxn_opcodes_h_l1045_c2_548e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1045_c2_548e_cond <= VAR_n8_MUX_uxn_opcodes_h_l1045_c2_548e_cond;
     n8_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue;
     n8_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1045_c2_548e_return_output := n8_MUX_uxn_opcodes_h_l1045_c2_548e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1045_c2_548e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1045_c2_548e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1050_c7_eab2_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1045_c2_548e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1045_c2_548e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1045_c2_548e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1074_l1041_DUPLICATE_34fe LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1074_l1041_DUPLICATE_34fe_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_641b(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1045_c2_548e_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1045_c2_548e_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1045_c2_548e_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1045_c2_548e_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1045_c2_548e_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1045_c2_548e_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1074_l1041_DUPLICATE_34fe_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1074_l1041_DUPLICATE_34fe_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
