-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity opc_sta_phased_0CLK_315c45c0 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(3 downto 0);
 pc : in unsigned(15 downto 0);
 sp : in unsigned(7 downto 0);
 stack_index : in unsigned(0 downto 0);
 ins : in unsigned(7 downto 0);
 k : in unsigned(7 downto 0);
 return_output : out unsigned(0 downto 0));
end opc_sta_phased_0CLK_315c45c0;
architecture arch of opc_sta_phased_0CLK_315c45c0 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal l8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal set_will_succeed : unsigned(0 downto 0) := to_unsigned(0, 1);
signal result : unsigned(0 downto 0) := to_unsigned(0, 1);
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_l8 : unsigned(7 downto 0);
signal REG_COMB_set_will_succeed : unsigned(0 downto 0);
signal REG_COMB_result : unsigned(0 downto 0);

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_phased_h_l833_c6_e73e]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l833_c1_ebb5]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l836_c7_ff51]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_phased_h_l833_c2_570d]
signal t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_return_output : unsigned(15 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l833_c2_570d]
signal result_MUX_uxn_opcodes_phased_h_l833_c2_570d_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l833_c2_570d_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l833_c2_570d_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l833_c2_570d_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_phased_h_l833_c2_570d]
signal l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_return_output : unsigned(7 downto 0);

-- set_will_fail[uxn_opcodes_phased_h_l834_c12_e535]
signal set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_sp : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_k : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_mul : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_add : signed(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l836_c11_6a74]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l836_c1_cfdc]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l839_c7_11dd]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_phased_h_l836_c7_ff51]
signal t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output : unsigned(15 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l836_c7_ff51]
signal result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_phased_h_l836_c7_ff51]
signal l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output : unsigned(7 downto 0);

-- t2_register[uxn_opcodes_phased_h_l837_c9_7a25]
signal t2_register_uxn_opcodes_phased_h_l837_c9_7a25_CLOCK_ENABLE : unsigned(0 downto 0);
signal t2_register_uxn_opcodes_phased_h_l837_c9_7a25_stack_index : unsigned(0 downto 0);
signal t2_register_uxn_opcodes_phased_h_l837_c9_7a25_stack_ptr : unsigned(7 downto 0);
signal t2_register_uxn_opcodes_phased_h_l837_c9_7a25_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l839_c11_cfea]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l839_c1_2a5e]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l842_c7_0849]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_phased_h_l839_c7_11dd]
signal t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output : unsigned(15 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l839_c7_11dd]
signal result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_phased_h_l839_c7_11dd]
signal l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output : unsigned(7 downto 0);

-- t2_register[uxn_opcodes_phased_h_l840_c9_79fd]
signal t2_register_uxn_opcodes_phased_h_l840_c9_79fd_CLOCK_ENABLE : unsigned(0 downto 0);
signal t2_register_uxn_opcodes_phased_h_l840_c9_79fd_stack_index : unsigned(0 downto 0);
signal t2_register_uxn_opcodes_phased_h_l840_c9_79fd_stack_ptr : unsigned(7 downto 0);
signal t2_register_uxn_opcodes_phased_h_l840_c9_79fd_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l842_c11_f79d]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l842_c11_f79d_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l842_c11_f79d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l842_c11_f79d_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l842_c1_daa8]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l845_c7_4ac0]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l842_c7_0849]
signal result_MUX_uxn_opcodes_phased_h_l842_c7_0849_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l842_c7_0849_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l842_c7_0849_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l842_c7_0849_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_phased_h_l842_c7_0849]
signal l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_return_output : unsigned(7 downto 0);

-- l_register[uxn_opcodes_phased_h_l843_c8_6f96]
signal l_register_uxn_opcodes_phased_h_l843_c8_6f96_CLOCK_ENABLE : unsigned(0 downto 0);
signal l_register_uxn_opcodes_phased_h_l843_c8_6f96_stack_index : unsigned(0 downto 0);
signal l_register_uxn_opcodes_phased_h_l843_c8_6f96_stack_ptr : unsigned(7 downto 0);
signal l_register_uxn_opcodes_phased_h_l843_c8_6f96_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l845_c11_ed2a]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l845_c11_ed2a_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l845_c11_ed2a_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l845_c11_ed2a_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l845_c1_274e]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l848_c7_e217]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l845_c7_4ac0]
signal result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_phased_h_l845_c7_4ac0]
signal l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_return_output : unsigned(7 downto 0);

-- l_register[uxn_opcodes_phased_h_l846_c8_5f53]
signal l_register_uxn_opcodes_phased_h_l846_c8_5f53_CLOCK_ENABLE : unsigned(0 downto 0);
signal l_register_uxn_opcodes_phased_h_l846_c8_5f53_stack_index : unsigned(0 downto 0);
signal l_register_uxn_opcodes_phased_h_l846_c8_5f53_stack_ptr : unsigned(7 downto 0);
signal l_register_uxn_opcodes_phased_h_l846_c8_5f53_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l848_c11_7fd0]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l848_c11_7fd0_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l848_c11_7fd0_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l848_c11_7fd0_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l848_c1_66ff]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l848_c7_e217]
signal result_MUX_uxn_opcodes_phased_h_l848_c7_e217_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l848_c7_e217_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l848_c7_e217_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l848_c7_e217_return_output : unsigned(0 downto 0);

-- set[uxn_opcodes_phased_h_l849_c3_e795]
signal set_uxn_opcodes_phased_h_l849_c3_e795_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l849_c3_e795_sp : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l849_c3_e795_stack_index : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l849_c3_e795_ins : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l849_c3_e795_k : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l849_c3_e795_mul : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l849_c3_e795_add : signed(7 downto 0);

-- poke_ram[uxn_opcodes_phased_h_l850_c3_82e7]
signal poke_ram_uxn_opcodes_phased_h_l850_c3_82e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal poke_ram_uxn_opcodes_phased_h_l850_c3_82e7_address : unsigned(15 downto 0);
signal poke_ram_uxn_opcodes_phased_h_l850_c3_82e7_value : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l852_c11_cb43]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l852_c11_cb43_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l852_c11_cb43_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l852_c11_cb43_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l852_c7_bb78]
signal result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_return_output : unsigned(0 downto 0);


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e
BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output);

-- t16_MUX_uxn_opcodes_phased_h_l833_c2_570d
t16_MUX_uxn_opcodes_phased_h_l833_c2_570d : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_cond,
t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_iftrue,
t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_iffalse,
t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_return_output);

-- result_MUX_uxn_opcodes_phased_h_l833_c2_570d
result_MUX_uxn_opcodes_phased_h_l833_c2_570d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l833_c2_570d_cond,
result_MUX_uxn_opcodes_phased_h_l833_c2_570d_iftrue,
result_MUX_uxn_opcodes_phased_h_l833_c2_570d_iffalse,
result_MUX_uxn_opcodes_phased_h_l833_c2_570d_return_output);

-- l8_MUX_uxn_opcodes_phased_h_l833_c2_570d
l8_MUX_uxn_opcodes_phased_h_l833_c2_570d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_cond,
l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_iftrue,
l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_iffalse,
l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_return_output);

-- set_will_fail_uxn_opcodes_phased_h_l834_c12_e535
set_will_fail_uxn_opcodes_phased_h_l834_c12_e535 : entity work.set_will_fail_0CLK_23eb2db7 port map (
clk,
set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_CLOCK_ENABLE,
set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_sp,
set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_k,
set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_mul,
set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_add,
set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74
BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74 : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output);

-- t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51
t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_cond,
t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iftrue,
t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iffalse,
t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output);

-- result_MUX_uxn_opcodes_phased_h_l836_c7_ff51
result_MUX_uxn_opcodes_phased_h_l836_c7_ff51 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_cond,
result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iftrue,
result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iffalse,
result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output);

-- l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51
l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_cond,
l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iftrue,
l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iffalse,
l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output);

-- t2_register_uxn_opcodes_phased_h_l837_c9_7a25
t2_register_uxn_opcodes_phased_h_l837_c9_7a25 : entity work.t2_register_0CLK_a2cd5ea9 port map (
clk,
t2_register_uxn_opcodes_phased_h_l837_c9_7a25_CLOCK_ENABLE,
t2_register_uxn_opcodes_phased_h_l837_c9_7a25_stack_index,
t2_register_uxn_opcodes_phased_h_l837_c9_7a25_stack_ptr,
t2_register_uxn_opcodes_phased_h_l837_c9_7a25_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea
BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_return_output);

-- t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd
t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_cond,
t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iftrue,
t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iffalse,
t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output);

-- result_MUX_uxn_opcodes_phased_h_l839_c7_11dd
result_MUX_uxn_opcodes_phased_h_l839_c7_11dd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_cond,
result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iftrue,
result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iffalse,
result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output);

-- l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd
l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_cond,
l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iftrue,
l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iffalse,
l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output);

-- t2_register_uxn_opcodes_phased_h_l840_c9_79fd
t2_register_uxn_opcodes_phased_h_l840_c9_79fd : entity work.t2_register_0CLK_a2cd5ea9 port map (
clk,
t2_register_uxn_opcodes_phased_h_l840_c9_79fd_CLOCK_ENABLE,
t2_register_uxn_opcodes_phased_h_l840_c9_79fd_stack_index,
t2_register_uxn_opcodes_phased_h_l840_c9_79fd_stack_ptr,
t2_register_uxn_opcodes_phased_h_l840_c9_79fd_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l842_c11_f79d
BIN_OP_EQ_uxn_opcodes_phased_h_l842_c11_f79d : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l842_c11_f79d_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l842_c11_f79d_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l842_c11_f79d_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_return_output);

-- result_MUX_uxn_opcodes_phased_h_l842_c7_0849
result_MUX_uxn_opcodes_phased_h_l842_c7_0849 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l842_c7_0849_cond,
result_MUX_uxn_opcodes_phased_h_l842_c7_0849_iftrue,
result_MUX_uxn_opcodes_phased_h_l842_c7_0849_iffalse,
result_MUX_uxn_opcodes_phased_h_l842_c7_0849_return_output);

-- l8_MUX_uxn_opcodes_phased_h_l842_c7_0849
l8_MUX_uxn_opcodes_phased_h_l842_c7_0849 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_cond,
l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_iftrue,
l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_iffalse,
l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_return_output);

-- l_register_uxn_opcodes_phased_h_l843_c8_6f96
l_register_uxn_opcodes_phased_h_l843_c8_6f96 : entity work.l_register_0CLK_621d5f60 port map (
clk,
l_register_uxn_opcodes_phased_h_l843_c8_6f96_CLOCK_ENABLE,
l_register_uxn_opcodes_phased_h_l843_c8_6f96_stack_index,
l_register_uxn_opcodes_phased_h_l843_c8_6f96_stack_ptr,
l_register_uxn_opcodes_phased_h_l843_c8_6f96_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l845_c11_ed2a
BIN_OP_EQ_uxn_opcodes_phased_h_l845_c11_ed2a : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l845_c11_ed2a_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l845_c11_ed2a_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l845_c11_ed2a_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_return_output);

-- result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0
result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_cond,
result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iftrue,
result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iffalse,
result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_return_output);

-- l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0
l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_cond,
l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iftrue,
l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iffalse,
l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_return_output);

-- l_register_uxn_opcodes_phased_h_l846_c8_5f53
l_register_uxn_opcodes_phased_h_l846_c8_5f53 : entity work.l_register_0CLK_621d5f60 port map (
clk,
l_register_uxn_opcodes_phased_h_l846_c8_5f53_CLOCK_ENABLE,
l_register_uxn_opcodes_phased_h_l846_c8_5f53_stack_index,
l_register_uxn_opcodes_phased_h_l846_c8_5f53_stack_ptr,
l_register_uxn_opcodes_phased_h_l846_c8_5f53_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l848_c11_7fd0
BIN_OP_EQ_uxn_opcodes_phased_h_l848_c11_7fd0 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l848_c11_7fd0_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l848_c11_7fd0_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l848_c11_7fd0_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_return_output);

-- result_MUX_uxn_opcodes_phased_h_l848_c7_e217
result_MUX_uxn_opcodes_phased_h_l848_c7_e217 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l848_c7_e217_cond,
result_MUX_uxn_opcodes_phased_h_l848_c7_e217_iftrue,
result_MUX_uxn_opcodes_phased_h_l848_c7_e217_iffalse,
result_MUX_uxn_opcodes_phased_h_l848_c7_e217_return_output);

-- set_uxn_opcodes_phased_h_l849_c3_e795
set_uxn_opcodes_phased_h_l849_c3_e795 : entity work.set_0CLK_6f2c5aad port map (
clk,
set_uxn_opcodes_phased_h_l849_c3_e795_CLOCK_ENABLE,
set_uxn_opcodes_phased_h_l849_c3_e795_sp,
set_uxn_opcodes_phased_h_l849_c3_e795_stack_index,
set_uxn_opcodes_phased_h_l849_c3_e795_ins,
set_uxn_opcodes_phased_h_l849_c3_e795_k,
set_uxn_opcodes_phased_h_l849_c3_e795_mul,
set_uxn_opcodes_phased_h_l849_c3_e795_add);

-- poke_ram_uxn_opcodes_phased_h_l850_c3_82e7
poke_ram_uxn_opcodes_phased_h_l850_c3_82e7 : entity work.poke_ram_0CLK_de264c78 port map (
poke_ram_uxn_opcodes_phased_h_l850_c3_82e7_CLOCK_ENABLE,
poke_ram_uxn_opcodes_phased_h_l850_c3_82e7_address,
poke_ram_uxn_opcodes_phased_h_l850_c3_82e7_value);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l852_c11_cb43
BIN_OP_EQ_uxn_opcodes_phased_h_l852_c11_cb43 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l852_c11_cb43_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l852_c11_cb43_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l852_c11_cb43_return_output);

-- result_MUX_uxn_opcodes_phased_h_l852_c7_bb78
result_MUX_uxn_opcodes_phased_h_l852_c7_bb78 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_cond,
result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_iftrue,
result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_iffalse,
result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 sp,
 stack_index,
 ins,
 k,
 -- Registers
 t16,
 l8,
 set_will_succeed,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output,
 t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_return_output,
 result_MUX_uxn_opcodes_phased_h_l833_c2_570d_return_output,
 l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_return_output,
 set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output,
 t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output,
 result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output,
 l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output,
 t2_register_uxn_opcodes_phased_h_l837_c9_7a25_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_return_output,
 t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output,
 result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output,
 l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output,
 t2_register_uxn_opcodes_phased_h_l840_c9_79fd_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l842_c11_f79d_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_return_output,
 result_MUX_uxn_opcodes_phased_h_l842_c7_0849_return_output,
 l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_return_output,
 l_register_uxn_opcodes_phased_h_l843_c8_6f96_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l845_c11_ed2a_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_return_output,
 result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_return_output,
 l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_return_output,
 l_register_uxn_opcodes_phased_h_l846_c8_5f53_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l848_c11_7fd0_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_return_output,
 result_MUX_uxn_opcodes_phased_h_l848_c7_e217_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l852_c11_cb43_return_output,
 result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(0 downto 0);
 variable VAR_phase : unsigned(3 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_sp : unsigned(7 downto 0);
 variable VAR_stack_index : unsigned(0 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_k : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iffalse : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l833_c2_570d_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l833_c2_570d_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l833_c2_570d_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l833_c2_570d_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_cond : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_sp : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_k : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_mul : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_add : signed(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iffalse : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_cond : unsigned(0 downto 0);
 variable VAR_t2_register_uxn_opcodes_phased_h_l837_c9_7a25_stack_index : unsigned(0 downto 0);
 variable VAR_t2_register_uxn_opcodes_phased_h_l837_c9_7a25_stack_ptr : unsigned(7 downto 0);
 variable VAR_t2_register_uxn_opcodes_phased_h_l837_c9_7a25_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_t2_register_uxn_opcodes_phased_h_l837_c9_7a25_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_iffalse : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l842_c7_0849_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_cond : unsigned(0 downto 0);
 variable VAR_t2_register_uxn_opcodes_phased_h_l840_c9_79fd_stack_index : unsigned(0 downto 0);
 variable VAR_t2_register_uxn_opcodes_phased_h_l840_c9_79fd_stack_ptr : unsigned(7 downto 0);
 variable VAR_t2_register_uxn_opcodes_phased_h_l840_c9_79fd_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_t2_register_uxn_opcodes_phased_h_l840_c9_79fd_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l842_c11_f79d_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l842_c11_f79d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l842_c11_f79d_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l842_c7_0849_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l842_c7_0849_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l842_c7_0849_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_cond : unsigned(0 downto 0);
 variable VAR_l_register_uxn_opcodes_phased_h_l843_c8_6f96_stack_index : unsigned(0 downto 0);
 variable VAR_l_register_uxn_opcodes_phased_h_l843_c8_6f96_stack_ptr : unsigned(7 downto 0);
 variable VAR_l_register_uxn_opcodes_phased_h_l843_c8_6f96_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_l_register_uxn_opcodes_phased_h_l843_c8_6f96_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l845_c11_ed2a_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l845_c11_ed2a_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l845_c11_ed2a_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l848_c7_e217_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_cond : unsigned(0 downto 0);
 variable VAR_l_register_uxn_opcodes_phased_h_l846_c8_5f53_stack_index : unsigned(0 downto 0);
 variable VAR_l_register_uxn_opcodes_phased_h_l846_c8_5f53_stack_ptr : unsigned(7 downto 0);
 variable VAR_l_register_uxn_opcodes_phased_h_l846_c8_5f53_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_l_register_uxn_opcodes_phased_h_l846_c8_5f53_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l848_c11_7fd0_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l848_c11_7fd0_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l848_c11_7fd0_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l848_c7_e217_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l848_c7_e217_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l848_c7_e217_cond : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l849_c3_e795_sp : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l849_c3_e795_stack_index : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l849_c3_e795_ins : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l849_c3_e795_k : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l849_c3_e795_mul : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l849_c3_e795_add : signed(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l849_c3_e795_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_poke_ram_uxn_opcodes_phased_h_l850_c3_82e7_address : unsigned(15 downto 0);
 variable VAR_poke_ram_uxn_opcodes_phased_h_l850_c3_82e7_value : unsigned(7 downto 0);
 variable VAR_poke_ram_uxn_opcodes_phased_h_l850_c3_82e7_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l852_c11_cb43_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l852_c11_cb43_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l852_c11_cb43_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_cond : unsigned(0 downto 0);
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_l8 : unsigned(7 downto 0);
variable REG_VAR_set_will_succeed : unsigned(0 downto 0);
variable REG_VAR_result : unsigned(0 downto 0);
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_l8 := l8;
  REG_VAR_set_will_succeed := set_will_succeed;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_set_uxn_opcodes_phased_h_l849_c3_e795_mul := resize(to_unsigned(3, 2), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l848_c11_7fd0_right := to_unsigned(5, 3);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_iffalse := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74_right := to_unsigned(1, 1);
     VAR_set_uxn_opcodes_phased_h_l849_c3_e795_add := resize(to_signed(-3, 3), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l852_c11_cb43_right := to_unsigned(6, 3);
     VAR_result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_iftrue := to_unsigned(1, 1);
     VAR_set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_mul := resize(to_unsigned(3, 2), 8);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea_right := to_unsigned(2, 2);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_iffalse := to_unsigned(0, 1);
     VAR_set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_add := resize(to_signed(-3, 3), 8);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l845_c11_ed2a_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l842_c11_f79d_right := to_unsigned(3, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_sp := sp;
     VAR_stack_index := stack_index;
     VAR_ins := ins;
     VAR_k := k;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iffalse := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_iftrue := VAR_CLOCK_ENABLE;
     VAR_set_uxn_opcodes_phased_h_l849_c3_e795_ins := VAR_ins;
     VAR_set_uxn_opcodes_phased_h_l849_c3_e795_k := VAR_k;
     VAR_set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_k := VAR_k;
     VAR_l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iffalse := l8;
     VAR_poke_ram_uxn_opcodes_phased_h_l850_c3_82e7_value := l8;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l842_c11_f79d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l845_c11_ed2a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l848_c11_7fd0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l852_c11_cb43_left := VAR_phase;
     VAR_result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l842_c7_0849_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l848_c7_e217_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_iffalse := result;
     REG_VAR_set_will_succeed := set_will_succeed;
     VAR_l_register_uxn_opcodes_phased_h_l843_c8_6f96_stack_ptr := VAR_sp;
     VAR_l_register_uxn_opcodes_phased_h_l846_c8_5f53_stack_ptr := VAR_sp;
     VAR_set_uxn_opcodes_phased_h_l849_c3_e795_sp := VAR_sp;
     VAR_set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_sp := VAR_sp;
     VAR_t2_register_uxn_opcodes_phased_h_l837_c9_7a25_stack_ptr := VAR_sp;
     VAR_t2_register_uxn_opcodes_phased_h_l840_c9_79fd_stack_ptr := VAR_sp;
     VAR_l_register_uxn_opcodes_phased_h_l843_c8_6f96_stack_index := VAR_stack_index;
     VAR_l_register_uxn_opcodes_phased_h_l846_c8_5f53_stack_index := VAR_stack_index;
     VAR_set_uxn_opcodes_phased_h_l849_c3_e795_stack_index := VAR_stack_index;
     VAR_t2_register_uxn_opcodes_phased_h_l837_c9_7a25_stack_index := VAR_stack_index;
     VAR_t2_register_uxn_opcodes_phased_h_l840_c9_79fd_stack_index := VAR_stack_index;
     VAR_poke_ram_uxn_opcodes_phased_h_l850_c3_82e7_address := t16;
     VAR_t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iffalse := t16;
     -- BIN_OP_EQ[uxn_opcodes_phased_h_l839_c11_cfea] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l842_c11_f79d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l842_c11_f79d_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l842_c11_f79d_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l842_c11_f79d_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l842_c11_f79d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l842_c11_f79d_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l842_c11_f79d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l836_c11_6a74] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l852_c11_cb43] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l852_c11_cb43_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l852_c11_cb43_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l852_c11_cb43_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l852_c11_cb43_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l852_c11_cb43_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l852_c11_cb43_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l833_c6_e73e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l845_c11_ed2a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l845_c11_ed2a_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l845_c11_ed2a_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l845_c11_ed2a_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l845_c11_ed2a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l845_c11_ed2a_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l845_c11_ed2a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l848_c11_7fd0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l848_c11_7fd0_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l848_c11_7fd0_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l848_c11_7fd0_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l848_c11_7fd0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l848_c11_7fd0_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l848_c11_7fd0_return_output;

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e_return_output;
     VAR_l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l833_c2_570d_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e_return_output;
     VAR_t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l833_c6_e73e_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74_return_output;
     VAR_l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74_return_output;
     VAR_t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l836_c11_6a74_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea_return_output;
     VAR_l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea_return_output;
     VAR_t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l839_c11_cfea_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l842_c11_f79d_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l842_c11_f79d_return_output;
     VAR_l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l842_c11_f79d_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l842_c7_0849_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l842_c11_f79d_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l845_c11_ed2a_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l845_c11_ed2a_return_output;
     VAR_l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l845_c11_ed2a_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l845_c11_ed2a_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l848_c11_7fd0_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l848_c7_e217_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l848_c11_7fd0_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l852_c11_cb43_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l852_c7_bb78] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_cond;
     result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_iftrue;
     result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_return_output := result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l833_c1_ebb5] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l836_c7_ff51] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output;
     VAR_set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l833_c1_ebb5_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l848_c7_e217_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l852_c7_bb78_return_output;
     -- set_will_fail[uxn_opcodes_phased_h_l834_c12_e535] LATENCY=0
     -- Clock enable
     set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_CLOCK_ENABLE <= VAR_set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_CLOCK_ENABLE;
     -- Inputs
     set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_sp <= VAR_set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_sp;
     set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_k <= VAR_set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_k;
     set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_mul <= VAR_set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_mul;
     set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_add <= VAR_set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_add;
     -- Outputs
     VAR_set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_return_output := set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l848_c7_e217] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l848_c7_e217_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l848_c7_e217_cond;
     result_MUX_uxn_opcodes_phased_h_l848_c7_e217_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l848_c7_e217_iftrue;
     result_MUX_uxn_opcodes_phased_h_l848_c7_e217_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l848_c7_e217_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l848_c7_e217_return_output := result_MUX_uxn_opcodes_phased_h_l848_c7_e217_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l836_c1_cfdc] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l839_c7_11dd] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output;

     -- Submodule level 3
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output;
     VAR_t2_register_uxn_opcodes_phased_h_l837_c9_7a25_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l836_c1_cfdc_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l848_c7_e217_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l833_c2_570d_iftrue := VAR_set_will_fail_uxn_opcodes_phased_h_l834_c12_e535_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l842_c7_0849] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l845_c7_4ac0] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_cond;
     result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iftrue;
     result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_return_output := result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l839_c1_2a5e] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_return_output;

     -- t2_register[uxn_opcodes_phased_h_l837_c9_7a25] LATENCY=0
     -- Clock enable
     t2_register_uxn_opcodes_phased_h_l837_c9_7a25_CLOCK_ENABLE <= VAR_t2_register_uxn_opcodes_phased_h_l837_c9_7a25_CLOCK_ENABLE;
     -- Inputs
     t2_register_uxn_opcodes_phased_h_l837_c9_7a25_stack_index <= VAR_t2_register_uxn_opcodes_phased_h_l837_c9_7a25_stack_index;
     t2_register_uxn_opcodes_phased_h_l837_c9_7a25_stack_ptr <= VAR_t2_register_uxn_opcodes_phased_h_l837_c9_7a25_stack_ptr;
     -- Outputs
     VAR_t2_register_uxn_opcodes_phased_h_l837_c9_7a25_return_output := t2_register_uxn_opcodes_phased_h_l837_c9_7a25_return_output;

     -- Submodule level 4
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c7_0849_return_output;
     VAR_t2_register_uxn_opcodes_phased_h_l840_c9_79fd_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l839_c1_2a5e_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l842_c7_0849_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_return_output;
     VAR_t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iftrue := VAR_t2_register_uxn_opcodes_phased_h_l837_c9_7a25_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l842_c7_0849] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l842_c7_0849_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l842_c7_0849_cond;
     result_MUX_uxn_opcodes_phased_h_l842_c7_0849_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l842_c7_0849_iftrue;
     result_MUX_uxn_opcodes_phased_h_l842_c7_0849_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l842_c7_0849_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l842_c7_0849_return_output := result_MUX_uxn_opcodes_phased_h_l842_c7_0849_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l842_c1_daa8] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_return_output;

     -- t2_register[uxn_opcodes_phased_h_l840_c9_79fd] LATENCY=0
     -- Clock enable
     t2_register_uxn_opcodes_phased_h_l840_c9_79fd_CLOCK_ENABLE <= VAR_t2_register_uxn_opcodes_phased_h_l840_c9_79fd_CLOCK_ENABLE;
     -- Inputs
     t2_register_uxn_opcodes_phased_h_l840_c9_79fd_stack_index <= VAR_t2_register_uxn_opcodes_phased_h_l840_c9_79fd_stack_index;
     t2_register_uxn_opcodes_phased_h_l840_c9_79fd_stack_ptr <= VAR_t2_register_uxn_opcodes_phased_h_l840_c9_79fd_stack_ptr;
     -- Outputs
     VAR_t2_register_uxn_opcodes_phased_h_l840_c9_79fd_return_output := t2_register_uxn_opcodes_phased_h_l840_c9_79fd_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l845_c7_4ac0] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_return_output;

     -- Submodule level 5
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_return_output;
     VAR_l_register_uxn_opcodes_phased_h_l843_c8_6f96_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l842_c1_daa8_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l842_c7_0849_return_output;
     VAR_t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iftrue := VAR_t2_register_uxn_opcodes_phased_h_l840_c9_79fd_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l845_c1_274e] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_return_output;

     -- l_register[uxn_opcodes_phased_h_l843_c8_6f96] LATENCY=0
     -- Clock enable
     l_register_uxn_opcodes_phased_h_l843_c8_6f96_CLOCK_ENABLE <= VAR_l_register_uxn_opcodes_phased_h_l843_c8_6f96_CLOCK_ENABLE;
     -- Inputs
     l_register_uxn_opcodes_phased_h_l843_c8_6f96_stack_index <= VAR_l_register_uxn_opcodes_phased_h_l843_c8_6f96_stack_index;
     l_register_uxn_opcodes_phased_h_l843_c8_6f96_stack_ptr <= VAR_l_register_uxn_opcodes_phased_h_l843_c8_6f96_stack_ptr;
     -- Outputs
     VAR_l_register_uxn_opcodes_phased_h_l843_c8_6f96_return_output := l_register_uxn_opcodes_phased_h_l843_c8_6f96_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l848_c7_e217] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_return_output;

     -- t16_MUX[uxn_opcodes_phased_h_l839_c7_11dd] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_cond <= VAR_t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_cond;
     t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iftrue <= VAR_t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iftrue;
     t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iffalse <= VAR_t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output := t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l839_c7_11dd] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_cond;
     result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iftrue;
     result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output := result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output;

     -- Submodule level 6
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c7_e217_return_output;
     VAR_l_register_uxn_opcodes_phased_h_l846_c8_5f53_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l845_c1_274e_return_output;
     VAR_l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_iftrue := VAR_l_register_uxn_opcodes_phased_h_l843_c8_6f96_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output;
     VAR_t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iffalse := VAR_t16_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output;
     -- t16_MUX[uxn_opcodes_phased_h_l836_c7_ff51] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_cond <= VAR_t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_cond;
     t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iftrue <= VAR_t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iftrue;
     t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iffalse <= VAR_t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output := t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l836_c7_ff51] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_cond;
     result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iftrue;
     result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output := result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output;

     -- l_register[uxn_opcodes_phased_h_l846_c8_5f53] LATENCY=0
     -- Clock enable
     l_register_uxn_opcodes_phased_h_l846_c8_5f53_CLOCK_ENABLE <= VAR_l_register_uxn_opcodes_phased_h_l846_c8_5f53_CLOCK_ENABLE;
     -- Inputs
     l_register_uxn_opcodes_phased_h_l846_c8_5f53_stack_index <= VAR_l_register_uxn_opcodes_phased_h_l846_c8_5f53_stack_index;
     l_register_uxn_opcodes_phased_h_l846_c8_5f53_stack_ptr <= VAR_l_register_uxn_opcodes_phased_h_l846_c8_5f53_stack_ptr;
     -- Outputs
     VAR_l_register_uxn_opcodes_phased_h_l846_c8_5f53_return_output := l_register_uxn_opcodes_phased_h_l846_c8_5f53_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l848_c1_66ff] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_return_output;

     -- Submodule level 7
     VAR_poke_ram_uxn_opcodes_phased_h_l850_c3_82e7_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_return_output;
     VAR_set_uxn_opcodes_phased_h_l849_c3_e795_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l848_c1_66ff_return_output;
     VAR_l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iftrue := VAR_l_register_uxn_opcodes_phased_h_l846_c8_5f53_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l833_c2_570d_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output;
     VAR_t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_iffalse := VAR_t16_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output;
     -- set[uxn_opcodes_phased_h_l849_c3_e795] LATENCY=0
     -- Clock enable
     set_uxn_opcodes_phased_h_l849_c3_e795_CLOCK_ENABLE <= VAR_set_uxn_opcodes_phased_h_l849_c3_e795_CLOCK_ENABLE;
     -- Inputs
     set_uxn_opcodes_phased_h_l849_c3_e795_sp <= VAR_set_uxn_opcodes_phased_h_l849_c3_e795_sp;
     set_uxn_opcodes_phased_h_l849_c3_e795_stack_index <= VAR_set_uxn_opcodes_phased_h_l849_c3_e795_stack_index;
     set_uxn_opcodes_phased_h_l849_c3_e795_ins <= VAR_set_uxn_opcodes_phased_h_l849_c3_e795_ins;
     set_uxn_opcodes_phased_h_l849_c3_e795_k <= VAR_set_uxn_opcodes_phased_h_l849_c3_e795_k;
     set_uxn_opcodes_phased_h_l849_c3_e795_mul <= VAR_set_uxn_opcodes_phased_h_l849_c3_e795_mul;
     set_uxn_opcodes_phased_h_l849_c3_e795_add <= VAR_set_uxn_opcodes_phased_h_l849_c3_e795_add;
     -- Outputs

     -- result_MUX[uxn_opcodes_phased_h_l833_c2_570d] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l833_c2_570d_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l833_c2_570d_cond;
     result_MUX_uxn_opcodes_phased_h_l833_c2_570d_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l833_c2_570d_iftrue;
     result_MUX_uxn_opcodes_phased_h_l833_c2_570d_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l833_c2_570d_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l833_c2_570d_return_output := result_MUX_uxn_opcodes_phased_h_l833_c2_570d_return_output;

     -- poke_ram[uxn_opcodes_phased_h_l850_c3_82e7] LATENCY=0
     -- Clock enable
     poke_ram_uxn_opcodes_phased_h_l850_c3_82e7_CLOCK_ENABLE <= VAR_poke_ram_uxn_opcodes_phased_h_l850_c3_82e7_CLOCK_ENABLE;
     -- Inputs
     poke_ram_uxn_opcodes_phased_h_l850_c3_82e7_address <= VAR_poke_ram_uxn_opcodes_phased_h_l850_c3_82e7_address;
     poke_ram_uxn_opcodes_phased_h_l850_c3_82e7_value <= VAR_poke_ram_uxn_opcodes_phased_h_l850_c3_82e7_value;
     -- Outputs

     -- l8_MUX[uxn_opcodes_phased_h_l845_c7_4ac0] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_cond <= VAR_l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_cond;
     l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iftrue <= VAR_l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iftrue;
     l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iffalse <= VAR_l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_return_output := l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_return_output;

     -- t16_MUX[uxn_opcodes_phased_h_l833_c2_570d] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_cond <= VAR_t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_cond;
     t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_iftrue <= VAR_t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_iftrue;
     t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_iffalse <= VAR_t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_return_output := t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_return_output;

     -- Submodule level 8
     VAR_l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_iffalse := VAR_l8_MUX_uxn_opcodes_phased_h_l845_c7_4ac0_return_output;
     REG_VAR_result := VAR_result_MUX_uxn_opcodes_phased_h_l833_c2_570d_return_output;
     VAR_return_output := VAR_result_MUX_uxn_opcodes_phased_h_l833_c2_570d_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_phased_h_l833_c2_570d_return_output;
     -- l8_MUX[uxn_opcodes_phased_h_l842_c7_0849] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_cond <= VAR_l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_cond;
     l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_iftrue <= VAR_l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_iftrue;
     l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_iffalse <= VAR_l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_return_output := l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_return_output;

     -- Submodule level 9
     VAR_l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iffalse := VAR_l8_MUX_uxn_opcodes_phased_h_l842_c7_0849_return_output;
     -- l8_MUX[uxn_opcodes_phased_h_l839_c7_11dd] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_cond <= VAR_l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_cond;
     l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iftrue <= VAR_l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iftrue;
     l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iffalse <= VAR_l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output := l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output;

     -- Submodule level 10
     VAR_l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iffalse := VAR_l8_MUX_uxn_opcodes_phased_h_l839_c7_11dd_return_output;
     -- l8_MUX[uxn_opcodes_phased_h_l836_c7_ff51] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_cond <= VAR_l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_cond;
     l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iftrue <= VAR_l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iftrue;
     l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iffalse <= VAR_l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output := l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output;

     -- Submodule level 11
     VAR_l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_iffalse := VAR_l8_MUX_uxn_opcodes_phased_h_l836_c7_ff51_return_output;
     -- l8_MUX[uxn_opcodes_phased_h_l833_c2_570d] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_cond <= VAR_l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_cond;
     l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_iftrue <= VAR_l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_iftrue;
     l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_iffalse <= VAR_l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_return_output := l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_return_output;

     -- Submodule level 12
     REG_VAR_l8 := VAR_l8_MUX_uxn_opcodes_phased_h_l833_c2_570d_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_l8 <= REG_VAR_l8;
REG_COMB_set_will_succeed <= REG_VAR_set_will_succeed;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     l8 <= REG_COMB_l8;
     set_will_succeed <= REG_COMB_set_will_succeed;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
