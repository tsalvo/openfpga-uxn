-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 53
entity lth_0CLK_6d7675a8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end lth_0CLK_6d7675a8;
architecture arch of lth_0CLK_6d7675a8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2004_c6_2dbe]
signal BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2004_c1_1df6]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2004_c2_4685]
signal n8_MUX_uxn_opcodes_h_l2004_c2_4685_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2004_c2_4685_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2004_c2_4685]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2004_c2_4685]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2004_c2_4685]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2004_c2_4685]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2004_c2_4685]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2004_c2_4685]
signal result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2004_c2_4685]
signal t8_MUX_uxn_opcodes_h_l2004_c2_4685_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2004_c2_4685_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l2005_c3_d6a5[uxn_opcodes_h_l2005_c3_d6a5]
signal printf_uxn_opcodes_h_l2005_c3_d6a5_uxn_opcodes_h_l2005_c3_d6a5_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2009_c11_2721]
signal BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2009_c7_bca0]
signal n8_MUX_uxn_opcodes_h_l2009_c7_bca0_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2009_c7_bca0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2009_c7_bca0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2009_c7_bca0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2009_c7_bca0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2009_c7_bca0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2009_c7_bca0]
signal result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2009_c7_bca0]
signal t8_MUX_uxn_opcodes_h_l2009_c7_bca0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2012_c11_93e3]
signal BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2012_c7_cd87]
signal n8_MUX_uxn_opcodes_h_l2012_c7_cd87_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2012_c7_cd87]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2012_c7_cd87]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2012_c7_cd87]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2012_c7_cd87]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2012_c7_cd87]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2012_c7_cd87]
signal result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2012_c7_cd87]
signal t8_MUX_uxn_opcodes_h_l2012_c7_cd87_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2016_c11_65a8]
signal BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2016_c7_78f2]
signal n8_MUX_uxn_opcodes_h_l2016_c7_78f2_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2016_c7_78f2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2016_c7_78f2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2016_c7_78f2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2016_c7_78f2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2016_c7_78f2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2016_c7_78f2]
signal result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2019_c11_c315]
signal BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2019_c7_f894]
signal n8_MUX_uxn_opcodes_h_l2019_c7_f894_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2019_c7_f894_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2019_c7_f894]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2019_c7_f894]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2019_c7_f894]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2019_c7_f894]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2019_c7_f894]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2019_c7_f894]
signal result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2022_c30_d09f]
signal sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_return_output : signed(3 downto 0);

-- BIN_OP_LT[uxn_opcodes_h_l2025_c21_9ad6]
signal BIN_OP_LT_uxn_opcodes_h_l2025_c21_9ad6_left : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l2025_c21_9ad6_right : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l2025_c21_9ad6_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l2025_c21_7a1b]
signal MUX_uxn_opcodes_h_l2025_c21_7a1b_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l2025_c21_7a1b_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l2025_c21_7a1b_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l2025_c21_7a1b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2027_c11_6ad9]
signal BIN_OP_EQ_uxn_opcodes_h_l2027_c11_6ad9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2027_c11_6ad9_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2027_c11_6ad9_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2027_c7_4bca]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2027_c7_4bca]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2027_c7_4bca]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8cda( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe
BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_left,
BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_right,
BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_return_output);

-- n8_MUX_uxn_opcodes_h_l2004_c2_4685
n8_MUX_uxn_opcodes_h_l2004_c2_4685 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2004_c2_4685_cond,
n8_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue,
n8_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse,
n8_MUX_uxn_opcodes_h_l2004_c2_4685_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685
result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685
result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685
result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685
result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685
result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_cond,
result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_return_output);

-- t8_MUX_uxn_opcodes_h_l2004_c2_4685
t8_MUX_uxn_opcodes_h_l2004_c2_4685 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2004_c2_4685_cond,
t8_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue,
t8_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse,
t8_MUX_uxn_opcodes_h_l2004_c2_4685_return_output);

-- printf_uxn_opcodes_h_l2005_c3_d6a5_uxn_opcodes_h_l2005_c3_d6a5
printf_uxn_opcodes_h_l2005_c3_d6a5_uxn_opcodes_h_l2005_c3_d6a5 : entity work.printf_uxn_opcodes_h_l2005_c3_d6a5_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2005_c3_d6a5_uxn_opcodes_h_l2005_c3_d6a5_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721
BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_left,
BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_right,
BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_return_output);

-- n8_MUX_uxn_opcodes_h_l2009_c7_bca0
n8_MUX_uxn_opcodes_h_l2009_c7_bca0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2009_c7_bca0_cond,
n8_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue,
n8_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse,
n8_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0
result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0
result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0
result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0
result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0
result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_cond,
result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output);

-- t8_MUX_uxn_opcodes_h_l2009_c7_bca0
t8_MUX_uxn_opcodes_h_l2009_c7_bca0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2009_c7_bca0_cond,
t8_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue,
t8_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse,
t8_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3
BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_left,
BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_right,
BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_return_output);

-- n8_MUX_uxn_opcodes_h_l2012_c7_cd87
n8_MUX_uxn_opcodes_h_l2012_c7_cd87 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2012_c7_cd87_cond,
n8_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue,
n8_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse,
n8_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87
result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87
result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87
result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87
result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87
result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_cond,
result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output);

-- t8_MUX_uxn_opcodes_h_l2012_c7_cd87
t8_MUX_uxn_opcodes_h_l2012_c7_cd87 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2012_c7_cd87_cond,
t8_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue,
t8_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse,
t8_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8
BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_left,
BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_right,
BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_return_output);

-- n8_MUX_uxn_opcodes_h_l2016_c7_78f2
n8_MUX_uxn_opcodes_h_l2016_c7_78f2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2016_c7_78f2_cond,
n8_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue,
n8_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse,
n8_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2
result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2
result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2
result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2
result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2
result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_cond,
result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315
BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_left,
BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_right,
BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_return_output);

-- n8_MUX_uxn_opcodes_h_l2019_c7_f894
n8_MUX_uxn_opcodes_h_l2019_c7_f894 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2019_c7_f894_cond,
n8_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue,
n8_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse,
n8_MUX_uxn_opcodes_h_l2019_c7_f894_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894
result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894
result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894
result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894
result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894
result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_cond,
result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f
sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_ins,
sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_x,
sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_y,
sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_return_output);

-- BIN_OP_LT_uxn_opcodes_h_l2025_c21_9ad6
BIN_OP_LT_uxn_opcodes_h_l2025_c21_9ad6 : entity work.BIN_OP_LT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_LT_uxn_opcodes_h_l2025_c21_9ad6_left,
BIN_OP_LT_uxn_opcodes_h_l2025_c21_9ad6_right,
BIN_OP_LT_uxn_opcodes_h_l2025_c21_9ad6_return_output);

-- MUX_uxn_opcodes_h_l2025_c21_7a1b
MUX_uxn_opcodes_h_l2025_c21_7a1b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l2025_c21_7a1b_cond,
MUX_uxn_opcodes_h_l2025_c21_7a1b_iftrue,
MUX_uxn_opcodes_h_l2025_c21_7a1b_iffalse,
MUX_uxn_opcodes_h_l2025_c21_7a1b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2027_c11_6ad9
BIN_OP_EQ_uxn_opcodes_h_l2027_c11_6ad9 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2027_c11_6ad9_left,
BIN_OP_EQ_uxn_opcodes_h_l2027_c11_6ad9_right,
BIN_OP_EQ_uxn_opcodes_h_l2027_c11_6ad9_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca
result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca
result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca
result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_return_output,
 n8_MUX_uxn_opcodes_h_l2004_c2_4685_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_return_output,
 t8_MUX_uxn_opcodes_h_l2004_c2_4685_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_return_output,
 n8_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output,
 t8_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_return_output,
 n8_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output,
 t8_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_return_output,
 n8_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_return_output,
 n8_MUX_uxn_opcodes_h_l2019_c7_f894_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_return_output,
 sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_return_output,
 BIN_OP_LT_uxn_opcodes_h_l2025_c21_9ad6_return_output,
 MUX_uxn_opcodes_h_l2025_c21_7a1b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2027_c11_6ad9_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2004_c2_4685_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2004_c2_4685_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2006_c3_6ac1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2004_c2_4685_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2004_c2_4685_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2005_c3_d6a5_uxn_opcodes_h_l2005_c3_d6a5_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2009_c7_bca0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2010_c3_e640 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2009_c7_bca0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2012_c7_cd87_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2014_c3_344a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2012_c7_cd87_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2019_c7_f894_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2016_c7_78f2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2017_c3_2cf9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2019_c7_f894_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2024_c3_9aaf : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2019_c7_f894_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2025_c21_7a1b_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2025_c21_7a1b_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2025_c21_7a1b_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l2025_c21_9ad6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l2025_c21_9ad6_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l2025_c21_9ad6_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2025_c21_7a1b_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2027_c11_6ad9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2027_c11_6ad9_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2027_c11_6ad9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2019_l2016_DUPLICATE_830c_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2027_l2016_DUPLICATE_cab3_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2027_l2016_DUPLICATE_f9e6_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2019_l2016_DUPLICATE_a589_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2012_l2009_l2027_l2019_l2016_DUPLICATE_01a0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l2000_l2033_DUPLICATE_4c67_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2017_c3_2cf9 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2017_c3_2cf9;
     VAR_sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2027_c11_6ad9_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2014_c3_344a := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2014_c3_344a;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2006_c3_6ac1 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2006_c3_6ac1;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_right := to_unsigned(4, 3);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_right := to_unsigned(3, 2);
     VAR_MUX_uxn_opcodes_h_l2025_c21_7a1b_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2010_c3_e640 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2010_c3_e640;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l2025_c21_7a1b_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2024_c3_9aaf := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2024_c3_9aaf;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2027_c11_6ad9_left := VAR_phase;
     VAR_BIN_OP_LT_uxn_opcodes_h_l2025_c21_9ad6_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_LT_uxn_opcodes_h_l2025_c21_9ad6_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2016_c11_65a8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_left;
     BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_return_output := BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2027_c11_6ad9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2027_c11_6ad9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2027_c11_6ad9_left;
     BIN_OP_EQ_uxn_opcodes_h_l2027_c11_6ad9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2027_c11_6ad9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2027_c11_6ad9_return_output := BIN_OP_EQ_uxn_opcodes_h_l2027_c11_6ad9_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2012_l2009_l2027_l2019_l2016_DUPLICATE_01a0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2012_l2009_l2027_l2019_l2016_DUPLICATE_01a0_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2027_l2016_DUPLICATE_cab3 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2027_l2016_DUPLICATE_cab3_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2012_c11_93e3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_left;
     BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_return_output := BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2009_c11_2721] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_left;
     BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_return_output := BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2019_c11_c315] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_left;
     BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_return_output := BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2004_c6_2dbe] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_left;
     BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_return_output := BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_return_output;

     -- BIN_OP_LT[uxn_opcodes_h_l2025_c21_9ad6] LATENCY=0
     -- Inputs
     BIN_OP_LT_uxn_opcodes_h_l2025_c21_9ad6_left <= VAR_BIN_OP_LT_uxn_opcodes_h_l2025_c21_9ad6_left;
     BIN_OP_LT_uxn_opcodes_h_l2025_c21_9ad6_right <= VAR_BIN_OP_LT_uxn_opcodes_h_l2025_c21_9ad6_right;
     -- Outputs
     VAR_BIN_OP_LT_uxn_opcodes_h_l2025_c21_9ad6_return_output := BIN_OP_LT_uxn_opcodes_h_l2025_c21_9ad6_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2019_l2016_DUPLICATE_830c LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2019_l2016_DUPLICATE_830c_return_output := result.sp_relative_shift;

     -- sp_relative_shift[uxn_opcodes_h_l2022_c30_d09f] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_ins;
     sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_x;
     sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_return_output := sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2019_l2016_DUPLICATE_a589 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2019_l2016_DUPLICATE_a589_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2027_l2016_DUPLICATE_f9e6 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2027_l2016_DUPLICATE_f9e6_return_output := result.is_stack_write;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2019_c7_f894] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2019_c7_f894_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2004_c2_4685_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2004_c2_4685_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2004_c6_2dbe_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2009_c7_bca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2009_c7_bca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c11_2721_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2012_c7_cd87_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2012_c7_cd87_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_93e3_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2016_c7_78f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2016_c11_65a8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2019_c7_f894_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_c315_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2027_c11_6ad9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2027_c11_6ad9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2027_c11_6ad9_return_output;
     VAR_MUX_uxn_opcodes_h_l2025_c21_7a1b_cond := VAR_BIN_OP_LT_uxn_opcodes_h_l2025_c21_9ad6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2019_l2016_DUPLICATE_830c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2019_l2016_DUPLICATE_830c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2019_l2016_DUPLICATE_830c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2019_l2016_DUPLICATE_830c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2019_l2016_DUPLICATE_830c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2012_l2009_l2027_l2019_l2016_DUPLICATE_01a0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2012_l2009_l2027_l2019_l2016_DUPLICATE_01a0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2012_l2009_l2027_l2019_l2016_DUPLICATE_01a0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2012_l2009_l2027_l2019_l2016_DUPLICATE_01a0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2012_l2009_l2027_l2019_l2016_DUPLICATE_01a0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2027_l2016_DUPLICATE_cab3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2027_l2016_DUPLICATE_cab3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2027_l2016_DUPLICATE_cab3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2027_l2016_DUPLICATE_cab3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2027_l2016_DUPLICATE_cab3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2027_l2016_DUPLICATE_f9e6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2027_l2016_DUPLICATE_f9e6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2027_l2016_DUPLICATE_f9e6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2027_l2016_DUPLICATE_f9e6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2027_l2016_DUPLICATE_f9e6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2019_l2016_DUPLICATE_a589_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2019_l2016_DUPLICATE_a589_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2019_l2016_DUPLICATE_a589_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2019_l2016_DUPLICATE_a589_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2012_l2009_l2004_l2019_l2016_DUPLICATE_a589_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2019_c7_f894_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2022_c30_d09f_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2027_c7_4bca] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2027_c7_4bca] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_return_output;

     -- MUX[uxn_opcodes_h_l2025_c21_7a1b] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l2025_c21_7a1b_cond <= VAR_MUX_uxn_opcodes_h_l2025_c21_7a1b_cond;
     MUX_uxn_opcodes_h_l2025_c21_7a1b_iftrue <= VAR_MUX_uxn_opcodes_h_l2025_c21_7a1b_iftrue;
     MUX_uxn_opcodes_h_l2025_c21_7a1b_iffalse <= VAR_MUX_uxn_opcodes_h_l2025_c21_7a1b_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l2025_c21_7a1b_return_output := MUX_uxn_opcodes_h_l2025_c21_7a1b_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2004_c1_1df6] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2019_c7_f894] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_return_output;

     -- t8_MUX[uxn_opcodes_h_l2012_c7_cd87] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2012_c7_cd87_cond <= VAR_t8_MUX_uxn_opcodes_h_l2012_c7_cd87_cond;
     t8_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue;
     t8_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output := t8_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2027_c7_4bca] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_return_output;

     -- n8_MUX[uxn_opcodes_h_l2019_c7_f894] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2019_c7_f894_cond <= VAR_n8_MUX_uxn_opcodes_h_l2019_c7_f894_cond;
     n8_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue;
     n8_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2019_c7_f894_return_output := n8_MUX_uxn_opcodes_h_l2019_c7_f894_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2019_c7_f894] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue := VAR_MUX_uxn_opcodes_h_l2025_c21_7a1b_return_output;
     VAR_printf_uxn_opcodes_h_l2005_c3_d6a5_uxn_opcodes_h_l2005_c3_d6a5_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2004_c1_1df6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2019_c7_f894_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2027_c7_4bca_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2027_c7_4bca_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2027_c7_4bca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_f894_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_f894_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2019_c7_f894] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_return_output;

     -- n8_MUX[uxn_opcodes_h_l2016_c7_78f2] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2016_c7_78f2_cond <= VAR_n8_MUX_uxn_opcodes_h_l2016_c7_78f2_cond;
     n8_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue;
     n8_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output := n8_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output;

     -- t8_MUX[uxn_opcodes_h_l2009_c7_bca0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2009_c7_bca0_cond <= VAR_t8_MUX_uxn_opcodes_h_l2009_c7_bca0_cond;
     t8_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue;
     t8_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output := t8_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2016_c7_78f2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2019_c7_f894] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_return_output;

     -- printf_uxn_opcodes_h_l2005_c3_d6a5[uxn_opcodes_h_l2005_c3_d6a5] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2005_c3_d6a5_uxn_opcodes_h_l2005_c3_d6a5_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2005_c3_d6a5_uxn_opcodes_h_l2005_c3_d6a5_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_u8_value_MUX[uxn_opcodes_h_l2019_c7_f894] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_return_output := result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2016_c7_78f2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2019_c7_f894] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_f894_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_f894_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_f894_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2019_c7_f894_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output;
     -- t8_MUX[uxn_opcodes_h_l2004_c2_4685] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2004_c2_4685_cond <= VAR_t8_MUX_uxn_opcodes_h_l2004_c2_4685_cond;
     t8_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue;
     t8_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2004_c2_4685_return_output := t8_MUX_uxn_opcodes_h_l2004_c2_4685_return_output;

     -- n8_MUX[uxn_opcodes_h_l2012_c7_cd87] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2012_c7_cd87_cond <= VAR_n8_MUX_uxn_opcodes_h_l2012_c7_cd87_cond;
     n8_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue;
     n8_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output := n8_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2016_c7_78f2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2012_c7_cd87] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2016_c7_78f2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output := result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2016_c7_78f2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2016_c7_78f2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2012_c7_cd87] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2016_c7_78f2_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2004_c2_4685_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2009_c7_bca0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2012_c7_cd87] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2012_c7_cd87] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2012_c7_cd87] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2012_c7_cd87] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output := result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output;

     -- n8_MUX[uxn_opcodes_h_l2009_c7_bca0] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2009_c7_bca0_cond <= VAR_n8_MUX_uxn_opcodes_h_l2009_c7_bca0_cond;
     n8_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue;
     n8_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output := n8_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2009_c7_bca0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2012_c7_cd87_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2009_c7_bca0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output := result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2009_c7_bca0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2009_c7_bca0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2004_c2_4685] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_return_output;

     -- n8_MUX[uxn_opcodes_h_l2004_c2_4685] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2004_c2_4685_cond <= VAR_n8_MUX_uxn_opcodes_h_l2004_c2_4685_cond;
     n8_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue;
     n8_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2004_c2_4685_return_output := n8_MUX_uxn_opcodes_h_l2004_c2_4685_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2009_c7_bca0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2004_c2_4685] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2004_c2_4685_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2009_c7_bca0_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2004_c2_4685] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2004_c2_4685] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2004_c2_4685] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2004_c2_4685] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_return_output := result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l2000_l2033_DUPLICATE_4c67 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l2000_l2033_DUPLICATE_4c67_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8cda(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2004_c2_4685_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2004_c2_4685_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2004_c2_4685_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2004_c2_4685_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2004_c2_4685_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2004_c2_4685_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l2000_l2033_DUPLICATE_4c67_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l2000_l2033_DUPLICATE_4c67_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
