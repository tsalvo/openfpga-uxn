-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 46
entity jsr_0CLK_fedec265 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jsr_0CLK_fedec265;
architecture arch of jsr_0CLK_fedec265 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l733_c6_2760]
signal BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l733_c2_9761]
signal result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l733_c2_9761]
signal result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l733_c2_9761]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_return_output : unsigned(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l733_c2_9761]
signal result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l733_c2_9761]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l733_c2_9761]
signal result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l733_c2_9761]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l733_c2_9761]
signal result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l733_c2_9761]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l733_c2_9761]
signal result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l733_c2_9761]
signal t8_MUX_uxn_opcodes_h_l733_c2_9761_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l733_c2_9761_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l733_c2_9761_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l733_c2_9761_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l746_c11_8a06]
signal BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l746_c7_6117]
signal result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l746_c7_6117]
signal result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l746_c7_6117]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l746_c7_6117]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_return_output : unsigned(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l746_c7_6117]
signal result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l746_c7_6117]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l746_c7_6117]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l746_c7_6117]
signal result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l746_c7_6117]
signal t8_MUX_uxn_opcodes_h_l746_c7_6117_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l746_c7_6117_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l746_c7_6117_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l746_c7_6117_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l748_c30_7586]
signal sp_relative_shift_uxn_opcodes_h_l748_c30_7586_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l748_c30_7586_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l748_c30_7586_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l748_c30_7586_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l750_c11_850c]
signal BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l750_c7_611f]
signal result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l750_c7_611f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l750_c7_611f]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l750_c7_611f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_return_output : unsigned(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l750_c7_611f]
signal result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l750_c7_611f]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l750_c7_611f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l750_c7_611f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l750_c7_611f]
signal t8_MUX_uxn_opcodes_h_l750_c7_611f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l750_c7_611f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l750_c7_611f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l750_c7_611f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l758_c11_9b6b]
signal BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l758_c7_5509]
signal result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l758_c7_5509]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_return_output : unsigned(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l758_c7_5509]
signal result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l758_c7_5509]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l758_c7_5509]
signal result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l758_c7_5509]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_return_output : unsigned(0 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l761_c31_0fb8]
signal CONST_SR_8_uxn_opcodes_h_l761_c31_0fb8_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l761_c31_0fb8_return_output : unsigned(15 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l763_c22_3e3d]
signal BIN_OP_PLUS_uxn_opcodes_h_l763_c22_3e3d_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l763_c22_3e3d_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l763_c22_3e3d_return_output : signed(17 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_2c6d( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : signed;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_vram_write := ref_toks_4;
      base.is_stack_index_flipped := ref_toks_5;
      base.u16_value := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.sp_relative_shift := ref_toks_9;
      base.is_opc_done := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760
BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_left,
BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_right,
BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761
result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_cond,
result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761
result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761
result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761
result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_cond,
result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761
result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761
result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761
result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761
result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_return_output);

-- t8_MUX_uxn_opcodes_h_l733_c2_9761
t8_MUX_uxn_opcodes_h_l733_c2_9761 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l733_c2_9761_cond,
t8_MUX_uxn_opcodes_h_l733_c2_9761_iftrue,
t8_MUX_uxn_opcodes_h_l733_c2_9761_iffalse,
t8_MUX_uxn_opcodes_h_l733_c2_9761_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06
BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_left,
BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_right,
BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117
result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_cond,
result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117
result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117
result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_cond,
result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117
result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117
result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117
result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_return_output);

-- t8_MUX_uxn_opcodes_h_l746_c7_6117
t8_MUX_uxn_opcodes_h_l746_c7_6117 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l746_c7_6117_cond,
t8_MUX_uxn_opcodes_h_l746_c7_6117_iftrue,
t8_MUX_uxn_opcodes_h_l746_c7_6117_iffalse,
t8_MUX_uxn_opcodes_h_l746_c7_6117_return_output);

-- sp_relative_shift_uxn_opcodes_h_l748_c30_7586
sp_relative_shift_uxn_opcodes_h_l748_c30_7586 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l748_c30_7586_ins,
sp_relative_shift_uxn_opcodes_h_l748_c30_7586_x,
sp_relative_shift_uxn_opcodes_h_l748_c30_7586_y,
sp_relative_shift_uxn_opcodes_h_l748_c30_7586_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c
BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_left,
BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_right,
BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f
result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_cond,
result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f
result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f
result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_cond,
result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f
result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f
result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f
result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_return_output);

-- t8_MUX_uxn_opcodes_h_l750_c7_611f
t8_MUX_uxn_opcodes_h_l750_c7_611f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l750_c7_611f_cond,
t8_MUX_uxn_opcodes_h_l750_c7_611f_iftrue,
t8_MUX_uxn_opcodes_h_l750_c7_611f_iffalse,
t8_MUX_uxn_opcodes_h_l750_c7_611f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b
BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b_left,
BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b_right,
BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509
result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_cond,
result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509
result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_cond,
result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509
result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509
result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509
result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_return_output);

-- CONST_SR_8_uxn_opcodes_h_l761_c31_0fb8
CONST_SR_8_uxn_opcodes_h_l761_c31_0fb8 : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l761_c31_0fb8_x,
CONST_SR_8_uxn_opcodes_h_l761_c31_0fb8_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l763_c22_3e3d
BIN_OP_PLUS_uxn_opcodes_h_l763_c22_3e3d : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l763_c22_3e3d_left,
BIN_OP_PLUS_uxn_opcodes_h_l763_c22_3e3d_right,
BIN_OP_PLUS_uxn_opcodes_h_l763_c22_3e3d_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_return_output,
 t8_MUX_uxn_opcodes_h_l733_c2_9761_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_return_output,
 t8_MUX_uxn_opcodes_h_l746_c7_6117_return_output,
 sp_relative_shift_uxn_opcodes_h_l748_c30_7586_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_return_output,
 t8_MUX_uxn_opcodes_h_l750_c7_611f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_return_output,
 CONST_SR_8_uxn_opcodes_h_l761_c31_0fb8_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l763_c22_3e3d_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l743_c3_3df7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l733_c2_9761_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l733_c2_9761_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l738_c3_80e6 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l733_c2_9761_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l733_c2_9761_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l746_c7_6117_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l733_c2_9761_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l733_c2_9761_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l747_c3_a059 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l746_c7_6117_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l746_c7_6117_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l750_c7_611f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l746_c7_6117_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l748_c30_7586_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l748_c30_7586_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l748_c30_7586_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l748_c30_7586_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l755_c3_d0bd : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l753_c3_43c2 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l750_c7_611f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l750_c7_611f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l750_c7_611f_cond : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l756_c21_5140_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l760_c3_0171 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l758_c7_5509_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l763_c3_0206 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l759_c3_44a4 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l758_c7_5509_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l761_c31_0fb8_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l761_c31_0fb8_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l761_c21_e810_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l763_c22_3e3d_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l763_c27_fd2c_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l763_c22_3e3d_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l763_c22_3e3d_return_output : signed(17 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l733_l758_l746_DUPLICATE_0f8e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l750_l733_l758_l746_DUPLICATE_ed6c_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l750_l746_DUPLICATE_1ece_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l750_l746_DUPLICATE_870a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l750_l758_l746_DUPLICATE_9895_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l750_l758_l746_DUPLICATE_7dd2_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_2c6d_uxn_opcodes_h_l767_l729_DUPLICATE_dc36_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l743_c3_3df7 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l743_c3_3df7;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l748_c30_7586_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l760_c3_0171 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l760_c3_0171;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l759_c3_44a4 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l759_c3_44a4;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l748_c30_7586_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l755_c3_d0bd := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l755_c3_d0bd;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_right := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_iftrue := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_right := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l738_c3_80e6 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l738_c3_80e6;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l753_c3_43c2 := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l753_c3_43c2;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l747_c3_a059 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l747_c3_a059;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l748_c30_7586_ins := VAR_ins;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l763_c22_3e3d_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_CONST_SR_8_uxn_opcodes_h_l761_c31_0fb8_x := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l750_c7_611f_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l733_c2_9761_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l746_c7_6117_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l750_c7_611f_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l750_l746_DUPLICATE_870a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l750_l746_DUPLICATE_870a_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l750_l746_DUPLICATE_1ece LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l750_l746_DUPLICATE_1ece_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l758_c11_9b6b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b_left;
     BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b_return_output := BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l733_l758_l746_DUPLICATE_0f8e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l733_l758_l746_DUPLICATE_0f8e_return_output := result.u8_value;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l758_c7_5509] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l758_c7_5509_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l733_c6_2760] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_left;
     BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_return_output := BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l733_c2_9761] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l733_c2_9761_return_output := result.is_ram_write;

     -- CONST_SR_8[uxn_opcodes_h_l761_c31_0fb8] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l761_c31_0fb8_x <= VAR_CONST_SR_8_uxn_opcodes_h_l761_c31_0fb8_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l761_c31_0fb8_return_output := CONST_SR_8_uxn_opcodes_h_l761_c31_0fb8_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l733_c2_9761] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l733_c2_9761_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l750_l758_l746_DUPLICATE_9895 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l750_l758_l746_DUPLICATE_9895_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l750_c11_850c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_left;
     BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_return_output := BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l746_c11_8a06] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_left;
     BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_return_output := BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_return_output;

     -- CAST_TO_int8_t[uxn_opcodes_h_l763_c27_fd2c] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l763_c27_fd2c_return_output := CAST_TO_int8_t_uint8_t(
     t8);

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l750_l758_l746_DUPLICATE_7dd2 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l750_l758_l746_DUPLICATE_7dd2_return_output := result.is_opc_done;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l756_c21_5140] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l756_c21_5140_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_pc);

     -- result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d[uxn_opcodes_h_l758_c7_5509] LATENCY=0
     VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l758_c7_5509_return_output := result.sp_relative_shift;

     -- sp_relative_shift[uxn_opcodes_h_l748_c30_7586] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l748_c30_7586_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l748_c30_7586_ins;
     sp_relative_shift_uxn_opcodes_h_l748_c30_7586_x <= VAR_sp_relative_shift_uxn_opcodes_h_l748_c30_7586_x;
     sp_relative_shift_uxn_opcodes_h_l748_c30_7586_y <= VAR_sp_relative_shift_uxn_opcodes_h_l748_c30_7586_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l748_c30_7586_return_output := sp_relative_shift_uxn_opcodes_h_l748_c30_7586_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l750_l733_l758_l746_DUPLICATE_ed6c LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l750_l733_l758_l746_DUPLICATE_ed6c_return_output := result.u16_value;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l733_c2_9761_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_2760_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l746_c7_6117_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_8a06_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l750_c7_611f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_850c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_9b6b_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l763_c22_3e3d_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l763_c27_fd2c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l756_c21_5140_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l750_l733_l758_l746_DUPLICATE_ed6c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l750_l733_l758_l746_DUPLICATE_ed6c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l750_l733_l758_l746_DUPLICATE_ed6c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l750_l733_l758_l746_DUPLICATE_ed6c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l750_l758_l746_DUPLICATE_7dd2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l750_l758_l746_DUPLICATE_7dd2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l750_l758_l746_DUPLICATE_7dd2_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l750_l758_l746_DUPLICATE_9895_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l750_l758_l746_DUPLICATE_9895_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l750_l758_l746_DUPLICATE_9895_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l750_l746_DUPLICATE_870a_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l750_l746_DUPLICATE_870a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l750_l746_DUPLICATE_1ece_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l750_l746_DUPLICATE_1ece_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l733_l758_l746_DUPLICATE_0f8e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l733_l758_l746_DUPLICATE_0f8e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l733_l758_l746_DUPLICATE_0f8e_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l733_c2_9761_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l733_c2_9761_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_iffalse := VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l758_c7_5509_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l758_c7_5509_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l748_c30_7586_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l758_c7_5509] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l758_c7_5509] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_return_output;

     -- t8_MUX[uxn_opcodes_h_l750_c7_611f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l750_c7_611f_cond <= VAR_t8_MUX_uxn_opcodes_h_l750_c7_611f_cond;
     t8_MUX_uxn_opcodes_h_l750_c7_611f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l750_c7_611f_iftrue;
     t8_MUX_uxn_opcodes_h_l750_c7_611f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l750_c7_611f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l750_c7_611f_return_output := t8_MUX_uxn_opcodes_h_l750_c7_611f_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l733_c2_9761] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l733_c2_9761] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l758_c7_5509] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l763_c22_3e3d] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l763_c22_3e3d_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l763_c22_3e3d_left;
     BIN_OP_PLUS_uxn_opcodes_h_l763_c22_3e3d_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l763_c22_3e3d_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l763_c22_3e3d_return_output := BIN_OP_PLUS_uxn_opcodes_h_l763_c22_3e3d_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l750_c7_611f] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l750_c7_611f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l758_c7_5509] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l761_c21_e810] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l761_c21_e810_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l761_c31_0fb8_return_output);

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l763_c3_0206 := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l763_c22_3e3d_return_output)),16);
     VAR_result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l761_c21_e810_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5509_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5509_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_611f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_611f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5509_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5509_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l746_c7_6117_iffalse := VAR_t8_MUX_uxn_opcodes_h_l750_c7_611f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_iftrue := VAR_result_u16_value_uxn_opcodes_h_l763_c3_0206;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l750_c7_611f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l750_c7_611f] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l750_c7_611f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l758_c7_5509] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_cond;
     result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_return_output := result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l746_c7_6117] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l758_c7_5509] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_cond;
     result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_return_output := result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l746_c7_6117] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_return_output;

     -- t8_MUX[uxn_opcodes_h_l746_c7_6117] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l746_c7_6117_cond <= VAR_t8_MUX_uxn_opcodes_h_l746_c7_6117_cond;
     t8_MUX_uxn_opcodes_h_l746_c7_6117_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l746_c7_6117_iftrue;
     t8_MUX_uxn_opcodes_h_l746_c7_6117_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l746_c7_6117_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l746_c7_6117_return_output := t8_MUX_uxn_opcodes_h_l746_c7_6117_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l750_c7_611f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_611f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_611f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_6117_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_6117_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_611f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_611f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l758_c7_5509_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l758_c7_5509_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l733_c2_9761_iffalse := VAR_t8_MUX_uxn_opcodes_h_l746_c7_6117_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l746_c7_6117] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l746_c7_6117] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l746_c7_6117] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l733_c2_9761] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l733_c2_9761] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l746_c7_6117] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_return_output;

     -- t8_MUX[uxn_opcodes_h_l733_c2_9761] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l733_c2_9761_cond <= VAR_t8_MUX_uxn_opcodes_h_l733_c2_9761_cond;
     t8_MUX_uxn_opcodes_h_l733_c2_9761_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l733_c2_9761_iftrue;
     t8_MUX_uxn_opcodes_h_l733_c2_9761_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l733_c2_9761_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l733_c2_9761_return_output := t8_MUX_uxn_opcodes_h_l733_c2_9761_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l750_c7_611f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_return_output := result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l750_c7_611f] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_cond;
     result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_return_output := result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_6117_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_6117_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_6117_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_6117_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_611f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_611f_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l733_c2_9761_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l733_c2_9761] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l733_c2_9761] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l733_c2_9761] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l746_c7_6117] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_cond;
     result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_return_output := result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l733_c2_9761] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l746_c7_6117] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_cond;
     result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_return_output := result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_return_output;

     -- Submodule level 5
     VAR_result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l746_c7_6117_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l746_c7_6117_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l733_c2_9761] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_cond;
     result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_return_output := result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l733_c2_9761] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_cond;
     result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_return_output := result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_2c6d_uxn_opcodes_h_l767_l729_DUPLICATE_dc36 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_2c6d_uxn_opcodes_h_l767_l729_DUPLICATE_dc36_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_2c6d(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l733_c2_9761_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_9761_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_9761_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_9761_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_9761_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l733_c2_9761_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_9761_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_9761_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_9761_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_9761_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_2c6d_uxn_opcodes_h_l767_l729_DUPLICATE_dc36_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_2c6d_uxn_opcodes_h_l767_l729_DUPLICATE_dc36_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
