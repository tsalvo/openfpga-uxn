-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 49
entity dei_0CLK_99af4b2a is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 controller0_buttons : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_device_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dei_0CLK_99af4b2a;
architecture arch of dei_0CLK_99af4b2a is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal has_written_to_t : unsigned(0 downto 0) := to_unsigned(0, 1);
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal device_in_result : device_in_result_t := device_in_result_t_NULL;
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_has_written_to_t : unsigned(0 downto 0);
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_device_in_result : device_in_result_t;
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l403_c6_20ab]
signal BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l419_c7_24d7]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l403_c2_2038]
signal t8_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(7 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l403_c2_2038]
signal has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(0 downto 0);

-- device_in_result_MUX[uxn_opcodes_h_l403_c2_2038]
signal device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
signal device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_return_output : device_in_result_t;

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l403_c2_2038]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l403_c2_2038]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l403_c2_2038]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l403_c2_2038]
signal result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(0 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l403_c2_2038]
signal result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l403_c2_2038]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l403_c2_2038]
signal result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l403_c2_2038]
signal result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l403_c2_2038]
signal result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l403_c2_2038]
signal result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(7 downto 0);

-- result_is_device_ram_write_MUX[uxn_opcodes_h_l403_c2_2038]
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l419_c11_0559]
signal BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l422_c1_ca63]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l419_c7_24d7]
signal t8_MUX_uxn_opcodes_h_l419_c7_24d7_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l419_c7_24d7_return_output : unsigned(7 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l419_c7_24d7]
signal has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_return_output : unsigned(0 downto 0);

-- device_in_result_MUX[uxn_opcodes_h_l419_c7_24d7]
signal device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_cond : unsigned(0 downto 0);
signal device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_return_output : device_in_result_t;

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l419_c7_24d7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l419_c7_24d7]
signal result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l419_c7_24d7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_return_output : unsigned(0 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l419_c7_24d7]
signal result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l419_c7_24d7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l419_c7_24d7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l420_c30_5631]
signal sp_relative_shift_uxn_opcodes_h_l420_c30_5631_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l420_c30_5631_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l420_c30_5631_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l420_c30_5631_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l424_c9_cd0c]
signal BIN_OP_EQ_uxn_opcodes_h_l424_c9_cd0c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l424_c9_cd0c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l424_c9_cd0c_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l424_c9_4a30]
signal MUX_uxn_opcodes_h_l424_c9_4a30_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l424_c9_4a30_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l424_c9_4a30_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l424_c9_4a30_return_output : unsigned(7 downto 0);

-- UNARY_OP_NOT[uxn_opcodes_h_l425_c8_8cc3]
signal UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8cc3_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8cc3_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l425_c1_6a15]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_return_output : unsigned(0 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l425_c3_6d3a]
signal has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output : unsigned(0 downto 0);

-- device_in_result_MUX[uxn_opcodes_h_l425_c3_6d3a]
signal device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_cond : unsigned(0 downto 0);
signal device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output : device_in_result_t;

-- result_u8_value_MUX[uxn_opcodes_h_l425_c3_6d3a]
signal result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l425_c3_6d3a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output : unsigned(0 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l425_c3_6d3a]
signal result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l425_c3_6d3a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l425_c3_6d3a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output : unsigned(0 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_h_l426_c37_8eb0]
signal BIN_OP_MINUS_uxn_opcodes_h_l426_c37_8eb0_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l426_c37_8eb0_right : unsigned(1 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l426_c37_8eb0_return_output : unsigned(7 downto 0);

-- device_in[uxn_opcodes_h_l426_c23_dbb2]
signal device_in_uxn_opcodes_h_l426_c23_dbb2_CLOCK_ENABLE : unsigned(0 downto 0);
signal device_in_uxn_opcodes_h_l426_c23_dbb2_device_address : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l426_c23_dbb2_phase : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l426_c23_dbb2_controller0_buttons : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l426_c23_dbb2_previous_device_ram_read : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l426_c23_dbb2_return_output : device_in_result_t;

-- UNARY_OP_NOT[uxn_opcodes_h_l429_c9_6048]
signal UNARY_OP_NOT_uxn_opcodes_h_l429_c9_6048_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_uxn_opcodes_h_l429_c9_6048_return_output : unsigned(0 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l429_c4_be04]
signal has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l429_c4_be04]
signal result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l429_c4_be04]
signal result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l429_c4_be04]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l429_c4_be04]
signal result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_return_output : unsigned(0 downto 0);

function CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6( ref_toks_0 : device_in_result_t;
 ref_toks_1 : unsigned) return device_in_result_t is
 
  variable base : device_in_result_t; 
  variable return_output : device_in_result_t;
begin
      base := ref_toks_0;
      base.is_dei_done := ref_toks_1;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_fa88( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.device_ram_address := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;
      base.is_opc_done := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.is_vram_write := ref_toks_9;
      base.u8_value := ref_toks_10;
      base.is_device_ram_write := ref_toks_11;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab
BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_left,
BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_right,
BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_return_output);

-- t8_MUX_uxn_opcodes_h_l403_c2_2038
t8_MUX_uxn_opcodes_h_l403_c2_2038 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l403_c2_2038_cond,
t8_MUX_uxn_opcodes_h_l403_c2_2038_iftrue,
t8_MUX_uxn_opcodes_h_l403_c2_2038_iffalse,
t8_MUX_uxn_opcodes_h_l403_c2_2038_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_cond,
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_return_output);

-- device_in_result_MUX_uxn_opcodes_h_l403_c2_2038
device_in_result_MUX_uxn_opcodes_h_l403_c2_2038 : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_cond,
device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_iftrue,
device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_iffalse,
device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038
result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_cond,
result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_return_output);

-- result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_cond,
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_iftrue,
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_iffalse,
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559
BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_left,
BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_right,
BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_return_output);

-- t8_MUX_uxn_opcodes_h_l419_c7_24d7
t8_MUX_uxn_opcodes_h_l419_c7_24d7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l419_c7_24d7_cond,
t8_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue,
t8_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse,
t8_MUX_uxn_opcodes_h_l419_c7_24d7_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_cond,
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_return_output);

-- device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7
device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7 : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_cond,
device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue,
device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse,
device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7
result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_cond,
result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_return_output);

-- sp_relative_shift_uxn_opcodes_h_l420_c30_5631
sp_relative_shift_uxn_opcodes_h_l420_c30_5631 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l420_c30_5631_ins,
sp_relative_shift_uxn_opcodes_h_l420_c30_5631_x,
sp_relative_shift_uxn_opcodes_h_l420_c30_5631_y,
sp_relative_shift_uxn_opcodes_h_l420_c30_5631_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l424_c9_cd0c
BIN_OP_EQ_uxn_opcodes_h_l424_c9_cd0c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l424_c9_cd0c_left,
BIN_OP_EQ_uxn_opcodes_h_l424_c9_cd0c_right,
BIN_OP_EQ_uxn_opcodes_h_l424_c9_cd0c_return_output);

-- MUX_uxn_opcodes_h_l424_c9_4a30
MUX_uxn_opcodes_h_l424_c9_4a30 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l424_c9_4a30_cond,
MUX_uxn_opcodes_h_l424_c9_4a30_iftrue,
MUX_uxn_opcodes_h_l424_c9_4a30_iffalse,
MUX_uxn_opcodes_h_l424_c9_4a30_return_output);

-- UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8cc3
UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8cc3 : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8cc3_expr,
UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8cc3_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_cond,
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output);

-- device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a
device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_cond,
device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue,
device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse,
device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a
result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_cond,
result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l426_c37_8eb0
BIN_OP_MINUS_uxn_opcodes_h_l426_c37_8eb0 : entity work.BIN_OP_MINUS_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l426_c37_8eb0_left,
BIN_OP_MINUS_uxn_opcodes_h_l426_c37_8eb0_right,
BIN_OP_MINUS_uxn_opcodes_h_l426_c37_8eb0_return_output);

-- device_in_uxn_opcodes_h_l426_c23_dbb2
device_in_uxn_opcodes_h_l426_c23_dbb2 : entity work.device_in_0CLK_50065acf port map (
clk,
device_in_uxn_opcodes_h_l426_c23_dbb2_CLOCK_ENABLE,
device_in_uxn_opcodes_h_l426_c23_dbb2_device_address,
device_in_uxn_opcodes_h_l426_c23_dbb2_phase,
device_in_uxn_opcodes_h_l426_c23_dbb2_controller0_buttons,
device_in_uxn_opcodes_h_l426_c23_dbb2_previous_device_ram_read,
device_in_uxn_opcodes_h_l426_c23_dbb2_return_output);

-- UNARY_OP_NOT_uxn_opcodes_h_l429_c9_6048
UNARY_OP_NOT_uxn_opcodes_h_l429_c9_6048 : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_uxn_opcodes_h_l429_c9_6048_expr,
UNARY_OP_NOT_uxn_opcodes_h_l429_c9_6048_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_cond,
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04
result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_cond,
result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 controller0_buttons,
 previous_stack_read,
 previous_device_ram_read,
 -- Registers
 has_written_to_t,
 t8,
 device_in_result,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_return_output,
 t8_MUX_uxn_opcodes_h_l403_c2_2038_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_return_output,
 device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_return_output,
 result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_return_output,
 t8_MUX_uxn_opcodes_h_l419_c7_24d7_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_return_output,
 device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_return_output,
 sp_relative_shift_uxn_opcodes_h_l420_c30_5631_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l424_c9_cd0c_return_output,
 MUX_uxn_opcodes_h_l424_c9_4a30_return_output,
 UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8cc3_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output,
 device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l426_c37_8eb0_return_output,
 device_in_uxn_opcodes_h_l426_c23_dbb2_return_output,
 UNARY_OP_NOT_uxn_opcodes_h_l429_c9_6048_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_controller0_buttons : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l419_c7_24d7_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : device_in_result_t;
 variable VAR_device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6_uxn_opcodes_h_l403_c2_2038_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l408_c3_8702 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l414_c3_e593 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l419_c7_24d7_cond : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_cond : unsigned(0 downto 0);
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l423_c3_bc3d : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_5631_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_5631_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_5631_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_5631_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l424_c9_4a30_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_cd0c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_cd0c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_cd0c_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l424_c9_4a30_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l424_c9_4a30_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l424_c9_4a30_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d_uxn_opcodes_h_l425_c8_9e92_return_output : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8cc3_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8cc3_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_cond : unsigned(0 downto 0);
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_cond : unsigned(0 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_dbb2_device_address : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_dbb2_phase : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_dbb2_controller0_buttons : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_dbb2_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_8eb0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_8eb0_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_8eb0_return_output : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_dbb2_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_dbb2_return_output : device_in_result_t;
 variable VAR_CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d_uxn_opcodes_h_l427_c32_8969_return_output : unsigned(7 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_6048_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_6048_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l431_c5_d882 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d_uxn_opcodes_h_l432_c23_55c0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l403_l425_l419_DUPLICATE_17f9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l403_l429_l425_l419_DUPLICATE_8d2c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l425_l419_DUPLICATE_f17d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l429_l425_l419_DUPLICATE_0574_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l429_l425_l419_DUPLICATE_ebcc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_fa88_uxn_opcodes_h_l397_l441_DUPLICATE_0509_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_has_written_to_t : unsigned(0 downto 0);
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_device_in_result : device_in_result_t;
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_has_written_to_t := has_written_to_t;
  REG_VAR_t8 := t8;
  REG_VAR_device_in_result := device_in_result;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_sp_relative_shift_uxn_opcodes_h_l423_c3_bc3d := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse := VAR_result_sp_relative_shift_uxn_opcodes_h_l423_c3_bc3d;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_iffalse := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l408_c3_8702 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l408_c3_8702;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l414_c3_e593 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l414_c3_e593;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_5631_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_8eb0_right := to_unsigned(2, 2);
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_cd0c_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_5631_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l431_c5_d882 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l431_c5_d882;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_right := to_unsigned(1, 1);
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_iftrue := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_controller0_buttons := controller0_buttons;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_device_ram_read := previous_device_ram_read;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse := VAR_CLOCK_ENABLE;
     VAR_device_in_uxn_opcodes_h_l426_c23_dbb2_controller0_buttons := VAR_controller0_buttons;
     VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue := device_in_result;
     VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse := device_in_result;
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_6048_expr := has_written_to_t;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue := has_written_to_t;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue := has_written_to_t;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_iffalse := has_written_to_t;
     VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_5631_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_cd0c_left := VAR_phase;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_8eb0_left := VAR_phase;
     VAR_device_in_uxn_opcodes_h_l426_c23_dbb2_previous_device_ram_read := VAR_previous_device_ram_read;
     VAR_MUX_uxn_opcodes_h_l424_c9_4a30_iftrue := VAR_previous_stack_read;
     VAR_MUX_uxn_opcodes_h_l424_c9_4a30_iffalse := t8;
     VAR_t8_MUX_uxn_opcodes_h_l403_c2_2038_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l424_c9_cd0c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l424_c9_cd0c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_cd0c_left;
     BIN_OP_EQ_uxn_opcodes_h_l424_c9_cd0c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_cd0c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_cd0c_return_output := BIN_OP_EQ_uxn_opcodes_h_l424_c9_cd0c_return_output;

     -- CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d[uxn_opcodes_h_l425_c8_9e92] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d_uxn_opcodes_h_l425_c8_9e92_return_output := device_in_result.is_dei_done;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l403_c2_2038] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l403_c2_2038_return_output := result.is_vram_write;

     -- sp_relative_shift[uxn_opcodes_h_l420_c30_5631] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l420_c30_5631_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_5631_ins;
     sp_relative_shift_uxn_opcodes_h_l420_c30_5631_x <= VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_5631_x;
     sp_relative_shift_uxn_opcodes_h_l420_c30_5631_y <= VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_5631_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_5631_return_output := sp_relative_shift_uxn_opcodes_h_l420_c30_5631_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l403_l429_l425_l419_DUPLICATE_8d2c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l403_l429_l425_l419_DUPLICATE_8d2c_return_output := result.u8_value;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l429_l425_l419_DUPLICATE_0574 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l429_l425_l419_DUPLICATE_0574_return_output := result.stack_address_sp_offset;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l403_c2_2038] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l403_c2_2038_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l403_c6_20ab] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_left;
     BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_return_output := BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_return_output;

     -- CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d[uxn_opcodes_h_l432_c23_55c0] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d_uxn_opcodes_h_l432_c23_55c0_return_output := device_in_result.dei_value;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l403_c2_2038] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l403_c2_2038_return_output := result.is_stack_index_flipped;

     -- UNARY_OP_NOT[uxn_opcodes_h_l429_c9_6048] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_uxn_opcodes_h_l429_c9_6048_expr <= VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_6048_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_6048_return_output := UNARY_OP_NOT_uxn_opcodes_h_l429_c9_6048_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l403_c2_2038] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l403_c2_2038_return_output := result.is_ram_write;

     -- BIN_OP_MINUS[uxn_opcodes_h_l426_c37_8eb0] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l426_c37_8eb0_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_8eb0_left;
     BIN_OP_MINUS_uxn_opcodes_h_l426_c37_8eb0_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_8eb0_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_8eb0_return_output := BIN_OP_MINUS_uxn_opcodes_h_l426_c37_8eb0_return_output;

     -- result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d[uxn_opcodes_h_l403_c2_2038] LATENCY=0
     VAR_result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l403_c2_2038_return_output := result.is_device_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l429_l425_l419_DUPLICATE_ebcc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l429_l425_l419_DUPLICATE_ebcc_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l425_l419_DUPLICATE_f17d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l425_l419_DUPLICATE_f17d_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l403_l425_l419_DUPLICATE_17f9 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l403_l425_l419_DUPLICATE_17f9_return_output := result.device_ram_address;

     -- device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6[uxn_opcodes_h_l403_c2_2038] LATENCY=0
     VAR_device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6_uxn_opcodes_h_l403_c2_2038_return_output := CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6(
     device_in_result,
     to_unsigned(0, 1));

     -- BIN_OP_EQ[uxn_opcodes_h_l419_c11_0559] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_left;
     BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_return_output := BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_return_output;

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l403_c2_2038_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_20ab_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l419_c7_24d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_0559_return_output;
     VAR_MUX_uxn_opcodes_h_l424_c9_4a30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_cd0c_return_output;
     VAR_device_in_uxn_opcodes_h_l426_c23_dbb2_phase := VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_8eb0_return_output;
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8cc3_expr := VAR_CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d_uxn_opcodes_h_l425_c8_9e92_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l429_l425_l419_DUPLICATE_ebcc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l429_l425_l419_DUPLICATE_ebcc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l429_l425_l419_DUPLICATE_ebcc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l425_l419_DUPLICATE_f17d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l425_l419_DUPLICATE_f17d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l429_l425_l419_DUPLICATE_0574_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l429_l425_l419_DUPLICATE_0574_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l429_l425_l419_DUPLICATE_0574_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_iftrue := VAR_CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d_uxn_opcodes_h_l432_c23_55c0_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l403_l425_l419_DUPLICATE_17f9_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l403_l425_l419_DUPLICATE_17f9_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l403_l425_l419_DUPLICATE_17f9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l403_l429_l425_l419_DUPLICATE_8d2c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l403_l429_l425_l419_DUPLICATE_8d2c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l403_l429_l425_l419_DUPLICATE_8d2c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l403_l429_l425_l419_DUPLICATE_8d2c_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_6048_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_6048_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_6048_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_6048_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_6048_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_iftrue := VAR_device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6_uxn_opcodes_h_l403_c2_2038_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_iffalse := VAR_result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l403_c2_2038_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l403_c2_2038_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l403_c2_2038_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l403_c2_2038_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l403_c2_2038_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_5631_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l419_c7_24d7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l429_c4_be04] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l429_c4_be04] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_cond;
     result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_return_output := result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l429_c4_be04] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_return_output := has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l403_c2_2038] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l403_c2_2038] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l419_c7_24d7] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l429_c4_be04] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l403_c2_2038] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output;

     -- MUX[uxn_opcodes_h_l424_c9_4a30] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l424_c9_4a30_cond <= VAR_MUX_uxn_opcodes_h_l424_c9_4a30_cond;
     MUX_uxn_opcodes_h_l424_c9_4a30_iftrue <= VAR_MUX_uxn_opcodes_h_l424_c9_4a30_iftrue;
     MUX_uxn_opcodes_h_l424_c9_4a30_iffalse <= VAR_MUX_uxn_opcodes_h_l424_c9_4a30_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l424_c9_4a30_return_output := MUX_uxn_opcodes_h_l424_c9_4a30_return_output;

     -- UNARY_OP_NOT[uxn_opcodes_h_l425_c8_8cc3] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8cc3_expr <= VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8cc3_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8cc3_return_output := UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8cc3_return_output;

     -- result_is_device_ram_write_MUX[uxn_opcodes_h_l403_c2_2038] LATENCY=0
     -- Inputs
     result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_cond <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_cond;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_iftrue <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_iftrue;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_iffalse <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_iffalse;
     -- Outputs
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output := result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l429_c4_be04] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l403_c2_2038] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_24d7_return_output;
     VAR_device_in_uxn_opcodes_h_l426_c23_dbb2_device_address := VAR_MUX_uxn_opcodes_h_l424_c9_4a30_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse := VAR_MUX_uxn_opcodes_h_l424_c9_4a30_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8cc3_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8cc3_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8cc3_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8cc3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8cc3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8cc3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8cc3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8cc3_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse := VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_be04_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_be04_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_be04_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_24d7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_be04_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_be04_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l403_c2_2038] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l422_c1_ca63] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l425_c3_6d3a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l425_c3_6d3a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output := result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l425_c3_6d3a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output;

     -- t8_MUX[uxn_opcodes_h_l419_c7_24d7] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l419_c7_24d7_cond <= VAR_t8_MUX_uxn_opcodes_h_l419_c7_24d7_cond;
     t8_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue;
     t8_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l419_c7_24d7_return_output := t8_MUX_uxn_opcodes_h_l419_c7_24d7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l425_c3_6d3a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l425_c3_6d3a] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output := has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output;

     -- Submodule level 3
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_ca63_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse := VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l403_c2_2038_iffalse := VAR_t8_MUX_uxn_opcodes_h_l419_c7_24d7_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l419_c7_24d7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_return_output;

     -- t8_MUX[uxn_opcodes_h_l403_c2_2038] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l403_c2_2038_cond <= VAR_t8_MUX_uxn_opcodes_h_l403_c2_2038_cond;
     t8_MUX_uxn_opcodes_h_l403_c2_2038_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l403_c2_2038_iftrue;
     t8_MUX_uxn_opcodes_h_l403_c2_2038_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l403_c2_2038_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l403_c2_2038_return_output := t8_MUX_uxn_opcodes_h_l403_c2_2038_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l419_c7_24d7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l425_c1_6a15] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l419_c7_24d7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l419_c7_24d7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_return_output := result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l419_c7_24d7] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_return_output := has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_return_output;

     -- Submodule level 4
     VAR_device_in_uxn_opcodes_h_l426_c23_dbb2_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_6a15_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_iffalse := VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_24d7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_24d7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_24d7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_24d7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_24d7_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l403_c2_2038_return_output;
     -- has_written_to_t_MUX[uxn_opcodes_h_l403_c2_2038] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_return_output := has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l403_c2_2038] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_cond;
     result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_return_output := result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l403_c2_2038] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l403_c2_2038] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l403_c2_2038] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output;

     -- device_in[uxn_opcodes_h_l426_c23_dbb2] LATENCY=0
     -- Clock enable
     device_in_uxn_opcodes_h_l426_c23_dbb2_CLOCK_ENABLE <= VAR_device_in_uxn_opcodes_h_l426_c23_dbb2_CLOCK_ENABLE;
     -- Inputs
     device_in_uxn_opcodes_h_l426_c23_dbb2_device_address <= VAR_device_in_uxn_opcodes_h_l426_c23_dbb2_device_address;
     device_in_uxn_opcodes_h_l426_c23_dbb2_phase <= VAR_device_in_uxn_opcodes_h_l426_c23_dbb2_phase;
     device_in_uxn_opcodes_h_l426_c23_dbb2_controller0_buttons <= VAR_device_in_uxn_opcodes_h_l426_c23_dbb2_controller0_buttons;
     device_in_uxn_opcodes_h_l426_c23_dbb2_previous_device_ram_read <= VAR_device_in_uxn_opcodes_h_l426_c23_dbb2_previous_device_ram_read;
     -- Outputs
     VAR_device_in_uxn_opcodes_h_l426_c23_dbb2_return_output := device_in_uxn_opcodes_h_l426_c23_dbb2_return_output;

     -- Submodule level 5
     VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue := VAR_device_in_uxn_opcodes_h_l426_c23_dbb2_return_output;
     REG_VAR_has_written_to_t := VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_2038_return_output;
     -- CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d[uxn_opcodes_h_l427_c32_8969] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d_uxn_opcodes_h_l427_c32_8969_return_output := VAR_device_in_uxn_opcodes_h_l426_c23_dbb2_return_output.device_ram_address;

     -- device_in_result_MUX[uxn_opcodes_h_l425_c3_6d3a] LATENCY=0
     -- Inputs
     device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_cond <= VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_cond;
     device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue <= VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue;
     device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse <= VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse;
     -- Outputs
     VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output := device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output;

     -- Submodule level 6
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue := VAR_CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d_uxn_opcodes_h_l427_c32_8969_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse := VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output;
     -- device_in_result_MUX[uxn_opcodes_h_l419_c7_24d7] LATENCY=0
     -- Inputs
     device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_cond <= VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_cond;
     device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue <= VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue;
     device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse <= VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse;
     -- Outputs
     VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_return_output := device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_return_output;

     -- result_device_ram_address_MUX[uxn_opcodes_h_l425_c3_6d3a] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output;

     -- Submodule level 7
     VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_iffalse := VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_24d7_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_6d3a_return_output;
     -- result_device_ram_address_MUX[uxn_opcodes_h_l419_c7_24d7] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_return_output;

     -- device_in_result_MUX[uxn_opcodes_h_l403_c2_2038] LATENCY=0
     -- Inputs
     device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_cond <= VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_cond;
     device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_iftrue <= VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_iftrue;
     device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_iffalse <= VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_iffalse;
     -- Outputs
     VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_return_output := device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_return_output;

     -- Submodule level 8
     REG_VAR_device_in_result := VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_2038_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_24d7_return_output;
     -- result_device_ram_address_MUX[uxn_opcodes_h_l403_c2_2038] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_return_output;

     -- Submodule level 9
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_fa88_uxn_opcodes_h_l397_l441_DUPLICATE_0509 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_fa88_uxn_opcodes_h_l397_l441_DUPLICATE_0509_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_fa88(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_2038_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_2038_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_2038_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output,
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_2038_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_2038_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_2038_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_2038_return_output,
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_2038_return_output);

     -- Submodule level 10
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_fa88_uxn_opcodes_h_l397_l441_DUPLICATE_0509_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_fa88_uxn_opcodes_h_l397_l441_DUPLICATE_0509_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_has_written_to_t <= REG_VAR_has_written_to_t;
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_device_in_result <= REG_VAR_device_in_result;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     has_written_to_t <= REG_COMB_has_written_to_t;
     t8 <= REG_COMB_t8;
     device_in_result <= REG_COMB_device_in_result;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
