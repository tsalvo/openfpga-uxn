-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 50
entity jmp2_0CLK_be70b838 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jmp2_0CLK_be70b838;
architecture arch of jmp2_0CLK_be70b838 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l654_c6_ac11]
signal BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l654_c1_22fc]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l654_c2_91dc]
signal t16_MUX_uxn_opcodes_h_l654_c2_91dc_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l654_c2_91dc_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l654_c2_91dc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l654_c2_91dc]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l654_c2_91dc]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l654_c2_91dc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l654_c2_91dc]
signal result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l654_c2_91dc]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_return_output : signed(3 downto 0);

-- printf_uxn_opcodes_h_l655_c3_b4df[uxn_opcodes_h_l655_c3_b4df]
signal printf_uxn_opcodes_h_l655_c3_b4df_uxn_opcodes_h_l655_c3_b4df_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l659_c11_bdc9]
signal BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l659_c7_a2a1]
signal t16_MUX_uxn_opcodes_h_l659_c7_a2a1_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l659_c7_a2a1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l659_c7_a2a1]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l659_c7_a2a1]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l659_c7_a2a1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l659_c7_a2a1]
signal result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l659_c7_a2a1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l662_c11_746a]
signal BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l662_c7_1277]
signal t16_MUX_uxn_opcodes_h_l662_c7_1277_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l662_c7_1277_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l662_c7_1277_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l662_c7_1277_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l662_c7_1277]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l662_c7_1277]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l662_c7_1277]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l662_c7_1277]
signal result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l662_c7_1277]
signal result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l662_c7_1277]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_return_output : signed(3 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l664_c3_8795]
signal CONST_SL_8_uxn_opcodes_h_l664_c3_8795_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l664_c3_8795_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l667_c11_fcd8]
signal BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l667_c7_ac90]
signal t16_MUX_uxn_opcodes_h_l667_c7_ac90_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l667_c7_ac90_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l667_c7_ac90]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l667_c7_ac90]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l667_c7_ac90]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l667_c7_ac90]
signal result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l667_c7_ac90]
signal result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l667_c7_ac90]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l670_c11_aed3]
signal BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l670_c7_bb45]
signal t16_MUX_uxn_opcodes_h_l670_c7_bb45_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l670_c7_bb45_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l670_c7_bb45]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l670_c7_bb45]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l670_c7_bb45]
signal result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l670_c7_bb45]
signal result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l670_c7_bb45]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_return_output : signed(3 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l671_c3_fc92]
signal BIN_OP_OR_uxn_opcodes_h_l671_c3_fc92_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l671_c3_fc92_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l671_c3_fc92_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l673_c30_d768]
signal sp_relative_shift_uxn_opcodes_h_l673_c30_d768_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l673_c30_d768_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l673_c30_d768_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l673_c30_d768_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l677_c11_f50e]
signal BIN_OP_EQ_uxn_opcodes_h_l677_c11_f50e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l677_c11_f50e_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l677_c11_f50e_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l677_c7_9df5]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l677_c7_9df5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l677_c7_9df5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_return_output : unsigned(0 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_8040( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.u16_value := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11
BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_left,
BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_right,
BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_return_output);

-- t16_MUX_uxn_opcodes_h_l654_c2_91dc
t16_MUX_uxn_opcodes_h_l654_c2_91dc : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l654_c2_91dc_cond,
t16_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue,
t16_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse,
t16_MUX_uxn_opcodes_h_l654_c2_91dc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc
result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc
result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc
result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc
result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_cond,
result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc
result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_return_output);

-- printf_uxn_opcodes_h_l655_c3_b4df_uxn_opcodes_h_l655_c3_b4df
printf_uxn_opcodes_h_l655_c3_b4df_uxn_opcodes_h_l655_c3_b4df : entity work.printf_uxn_opcodes_h_l655_c3_b4df_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l655_c3_b4df_uxn_opcodes_h_l655_c3_b4df_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9
BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_left,
BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_right,
BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_return_output);

-- t16_MUX_uxn_opcodes_h_l659_c7_a2a1
t16_MUX_uxn_opcodes_h_l659_c7_a2a1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l659_c7_a2a1_cond,
t16_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue,
t16_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse,
t16_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1
result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1
result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1
result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1
result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_cond,
result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1
result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a
BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_left,
BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_right,
BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_return_output);

-- t16_MUX_uxn_opcodes_h_l662_c7_1277
t16_MUX_uxn_opcodes_h_l662_c7_1277 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l662_c7_1277_cond,
t16_MUX_uxn_opcodes_h_l662_c7_1277_iftrue,
t16_MUX_uxn_opcodes_h_l662_c7_1277_iffalse,
t16_MUX_uxn_opcodes_h_l662_c7_1277_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277
result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277
result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277
result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277
result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_cond,
result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277
result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_return_output);

-- CONST_SL_8_uxn_opcodes_h_l664_c3_8795
CONST_SL_8_uxn_opcodes_h_l664_c3_8795 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l664_c3_8795_x,
CONST_SL_8_uxn_opcodes_h_l664_c3_8795_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8
BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_left,
BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_right,
BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_return_output);

-- t16_MUX_uxn_opcodes_h_l667_c7_ac90
t16_MUX_uxn_opcodes_h_l667_c7_ac90 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l667_c7_ac90_cond,
t16_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue,
t16_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse,
t16_MUX_uxn_opcodes_h_l667_c7_ac90_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90
result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90
result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90
result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90
result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_cond,
result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90
result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3
BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3_left,
BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3_right,
BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3_return_output);

-- t16_MUX_uxn_opcodes_h_l670_c7_bb45
t16_MUX_uxn_opcodes_h_l670_c7_bb45 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l670_c7_bb45_cond,
t16_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue,
t16_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse,
t16_MUX_uxn_opcodes_h_l670_c7_bb45_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45
result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45
result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45
result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45
result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_cond,
result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45
result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l671_c3_fc92
BIN_OP_OR_uxn_opcodes_h_l671_c3_fc92 : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l671_c3_fc92_left,
BIN_OP_OR_uxn_opcodes_h_l671_c3_fc92_right,
BIN_OP_OR_uxn_opcodes_h_l671_c3_fc92_return_output);

-- sp_relative_shift_uxn_opcodes_h_l673_c30_d768
sp_relative_shift_uxn_opcodes_h_l673_c30_d768 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l673_c30_d768_ins,
sp_relative_shift_uxn_opcodes_h_l673_c30_d768_x,
sp_relative_shift_uxn_opcodes_h_l673_c30_d768_y,
sp_relative_shift_uxn_opcodes_h_l673_c30_d768_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l677_c11_f50e
BIN_OP_EQ_uxn_opcodes_h_l677_c11_f50e : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l677_c11_f50e_left,
BIN_OP_EQ_uxn_opcodes_h_l677_c11_f50e_right,
BIN_OP_EQ_uxn_opcodes_h_l677_c11_f50e_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5
result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5
result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5
result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_return_output,
 t16_MUX_uxn_opcodes_h_l654_c2_91dc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_return_output,
 t16_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_return_output,
 t16_MUX_uxn_opcodes_h_l662_c7_1277_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_return_output,
 CONST_SL_8_uxn_opcodes_h_l664_c3_8795_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_return_output,
 t16_MUX_uxn_opcodes_h_l667_c7_ac90_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3_return_output,
 t16_MUX_uxn_opcodes_h_l670_c7_bb45_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_return_output,
 BIN_OP_OR_uxn_opcodes_h_l671_c3_fc92_return_output,
 sp_relative_shift_uxn_opcodes_h_l673_c30_d768_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l677_c11_f50e_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_iffalse : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l654_c2_91dc_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l654_c2_91dc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l656_c3_a57c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l655_c3_b4df_uxn_opcodes_h_l655_c3_b4df_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l662_c7_1277_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l659_c7_a2a1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l660_c3_8769 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l662_c7_1277_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l662_c7_1277_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l667_c7_ac90_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l662_c7_1277_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l665_c3_a57a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l664_c3_8795_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l664_c3_8795_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l670_c7_bb45_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l667_c7_ac90_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l668_c3_b2fa : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l667_c7_ac90_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l670_c7_bb45_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l671_c3_fc92_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l671_c3_fc92_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l671_c3_fc92_return_output : unsigned(15 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l673_c30_d768_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l673_c30_d768_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l673_c30_d768_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l673_c30_d768_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l677_c11_f50e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l677_c11_f50e_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l677_c11_f50e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l662_l659_l654_l677_l667_DUPLICATE_1c01_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l662_l659_l654_l677_l667_DUPLICATE_ee3f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l662_l659_l654_l667_l670_DUPLICATE_c946_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l662_l659_l654_l667_l670_DUPLICATE_2a9e_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l662_l659_l677_l667_l670_DUPLICATE_a9f6_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l663_l671_DUPLICATE_3f4b_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8040_uxn_opcodes_h_l683_l650_DUPLICATE_a750_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_right := to_unsigned(3, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l677_c11_f50e_right := to_unsigned(5, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l668_c3_b2fa := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l668_c3_b2fa;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l656_c3_a57c := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l656_c3_a57c;
     VAR_sp_relative_shift_uxn_opcodes_h_l673_c30_d768_y := resize(to_signed(-2, 3), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l660_c3_8769 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l660_c3_8769;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l665_c3_a57a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l665_c3_a57a;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l673_c30_d768_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_right := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l673_c30_d768_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l677_c11_f50e_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l671_c3_fc92_left := t16;
     VAR_t16_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse := t16;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l662_l659_l654_l677_l667_DUPLICATE_1c01 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l662_l659_l654_l677_l667_DUPLICATE_1c01_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l670_c11_aed3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3_left;
     BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3_return_output := BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l677_c11_f50e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l677_c11_f50e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l677_c11_f50e_left;
     BIN_OP_EQ_uxn_opcodes_h_l677_c11_f50e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l677_c11_f50e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l677_c11_f50e_return_output := BIN_OP_EQ_uxn_opcodes_h_l677_c11_f50e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l667_c11_fcd8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_left;
     BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_return_output := BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l662_l659_l654_l677_l667_DUPLICATE_ee3f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l662_l659_l654_l677_l667_DUPLICATE_ee3f_return_output := result.is_sp_shift;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l663_l671_DUPLICATE_3f4b LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l663_l671_DUPLICATE_3f4b_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l662_l659_l677_l667_l670_DUPLICATE_a9f6 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l662_l659_l677_l667_l670_DUPLICATE_a9f6_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l654_c6_ac11] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_left;
     BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_return_output := BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l659_c11_bdc9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_left;
     BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_return_output := BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l673_c30_d768] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l673_c30_d768_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l673_c30_d768_ins;
     sp_relative_shift_uxn_opcodes_h_l673_c30_d768_x <= VAR_sp_relative_shift_uxn_opcodes_h_l673_c30_d768_x;
     sp_relative_shift_uxn_opcodes_h_l673_c30_d768_y <= VAR_sp_relative_shift_uxn_opcodes_h_l673_c30_d768_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l673_c30_d768_return_output := sp_relative_shift_uxn_opcodes_h_l673_c30_d768_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l662_l659_l654_l667_l670_DUPLICATE_2a9e LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l662_l659_l654_l667_l670_DUPLICATE_2a9e_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l662_l659_l654_l667_l670_DUPLICATE_c946 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l662_l659_l654_l667_l670_DUPLICATE_c946_return_output := result.u16_value;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l667_c7_ac90] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l667_c7_ac90_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l662_c11_746a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_left;
     BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_return_output := BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l654_c2_91dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l654_c6_ac11_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l659_c7_a2a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l659_c11_bdc9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l662_c7_1277_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l662_c11_746a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l667_c7_ac90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l667_c11_fcd8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l670_c7_bb45_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l670_c11_aed3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l677_c11_f50e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l677_c11_f50e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l677_c11_f50e_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l671_c3_fc92_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l663_l671_DUPLICATE_3f4b_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l664_c3_8795_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l663_l671_DUPLICATE_3f4b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l662_l659_l654_l667_l670_DUPLICATE_2a9e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l662_l659_l654_l667_l670_DUPLICATE_2a9e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l662_l659_l654_l667_l670_DUPLICATE_2a9e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l662_l659_l654_l667_l670_DUPLICATE_2a9e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l662_l659_l654_l667_l670_DUPLICATE_2a9e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l662_l659_l654_l667_l670_DUPLICATE_c946_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l662_l659_l654_l667_l670_DUPLICATE_c946_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l662_l659_l654_l667_l670_DUPLICATE_c946_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l662_l659_l654_l667_l670_DUPLICATE_c946_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l662_l659_l654_l667_l670_DUPLICATE_c946_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l662_l659_l677_l667_l670_DUPLICATE_a9f6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l662_l659_l677_l667_l670_DUPLICATE_a9f6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l662_l659_l677_l667_l670_DUPLICATE_a9f6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l662_l659_l677_l667_l670_DUPLICATE_a9f6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l662_l659_l677_l667_l670_DUPLICATE_a9f6_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l662_l659_l654_l677_l667_DUPLICATE_1c01_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l662_l659_l654_l677_l667_DUPLICATE_1c01_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l662_l659_l654_l677_l667_DUPLICATE_1c01_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l662_l659_l654_l677_l667_DUPLICATE_1c01_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l662_l659_l654_l677_l667_DUPLICATE_1c01_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l662_l659_l654_l677_l667_DUPLICATE_ee3f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l662_l659_l654_l677_l667_DUPLICATE_ee3f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l662_l659_l654_l677_l667_DUPLICATE_ee3f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l662_l659_l654_l677_l667_DUPLICATE_ee3f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l662_l659_l654_l677_l667_DUPLICATE_ee3f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l667_c7_ac90_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l673_c30_d768_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l654_c1_22fc] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l677_c7_9df5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l664_c3_8795] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l664_c3_8795_x <= VAR_CONST_SL_8_uxn_opcodes_h_l664_c3_8795_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l664_c3_8795_return_output := CONST_SL_8_uxn_opcodes_h_l664_c3_8795_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l677_c7_9df5] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l670_c7_bb45] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l671_c3_fc92] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l671_c3_fc92_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l671_c3_fc92_left;
     BIN_OP_OR_uxn_opcodes_h_l671_c3_fc92_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l671_c3_fc92_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l671_c3_fc92_return_output := BIN_OP_OR_uxn_opcodes_h_l671_c3_fc92_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l677_c7_9df5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l667_c7_ac90] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_return_output;

     -- Submodule level 2
     VAR_result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l671_c3_fc92_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l671_c3_fc92_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l662_c7_1277_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l664_c3_8795_return_output;
     VAR_printf_uxn_opcodes_h_l655_c3_b4df_uxn_opcodes_h_l655_c3_b4df_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l654_c1_22fc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l677_c7_9df5_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l677_c7_9df5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l677_c7_9df5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l670_c7_bb45_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l667_c7_ac90_return_output;
     -- printf_uxn_opcodes_h_l655_c3_b4df[uxn_opcodes_h_l655_c3_b4df] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l655_c3_b4df_uxn_opcodes_h_l655_c3_b4df_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l655_c3_b4df_uxn_opcodes_h_l655_c3_b4df_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l667_c7_ac90] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l670_c7_bb45] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l670_c7_bb45] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_return_output;

     -- t16_MUX[uxn_opcodes_h_l670_c7_bb45] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l670_c7_bb45_cond <= VAR_t16_MUX_uxn_opcodes_h_l670_c7_bb45_cond;
     t16_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue;
     t16_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l670_c7_bb45_return_output := t16_MUX_uxn_opcodes_h_l670_c7_bb45_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l662_c7_1277] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l670_c7_bb45] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l670_c7_bb45] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_cond;
     result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_return_output := result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l670_c7_bb45_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l670_c7_bb45_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l670_c7_bb45_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l667_c7_ac90_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l662_c7_1277_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l670_c7_bb45_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse := VAR_t16_MUX_uxn_opcodes_h_l670_c7_bb45_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l667_c7_ac90] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_cond;
     result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_return_output := result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l662_c7_1277] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l667_c7_ac90] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l667_c7_ac90] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_return_output;

     -- t16_MUX[uxn_opcodes_h_l667_c7_ac90] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l667_c7_ac90_cond <= VAR_t16_MUX_uxn_opcodes_h_l667_c7_ac90_cond;
     t16_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue;
     t16_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l667_c7_ac90_return_output := t16_MUX_uxn_opcodes_h_l667_c7_ac90_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l659_c7_a2a1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l667_c7_ac90] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l667_c7_ac90_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l667_c7_ac90_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l667_c7_ac90_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l662_c7_1277_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l667_c7_ac90_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l662_c7_1277_iffalse := VAR_t16_MUX_uxn_opcodes_h_l667_c7_ac90_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l662_c7_1277] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_cond;
     result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_return_output := result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l662_c7_1277] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l662_c7_1277] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_return_output;

     -- t16_MUX[uxn_opcodes_h_l662_c7_1277] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l662_c7_1277_cond <= VAR_t16_MUX_uxn_opcodes_h_l662_c7_1277_cond;
     t16_MUX_uxn_opcodes_h_l662_c7_1277_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l662_c7_1277_iftrue;
     t16_MUX_uxn_opcodes_h_l662_c7_1277_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l662_c7_1277_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l662_c7_1277_return_output := t16_MUX_uxn_opcodes_h_l662_c7_1277_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l659_c7_a2a1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l662_c7_1277] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l654_c2_91dc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l662_c7_1277_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l662_c7_1277_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l662_c7_1277_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l662_c7_1277_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse := VAR_t16_MUX_uxn_opcodes_h_l662_c7_1277_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l659_c7_a2a1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l659_c7_a2a1] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output;

     -- t16_MUX[uxn_opcodes_h_l659_c7_a2a1] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l659_c7_a2a1_cond <= VAR_t16_MUX_uxn_opcodes_h_l659_c7_a2a1_cond;
     t16_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue;
     t16_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output := t16_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l659_c7_a2a1] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l654_c2_91dc] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l659_c7_a2a1] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_cond;
     result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output := result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse := VAR_t16_MUX_uxn_opcodes_h_l659_c7_a2a1_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l654_c2_91dc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_return_output;

     -- t16_MUX[uxn_opcodes_h_l654_c2_91dc] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l654_c2_91dc_cond <= VAR_t16_MUX_uxn_opcodes_h_l654_c2_91dc_cond;
     t16_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue;
     t16_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l654_c2_91dc_return_output := t16_MUX_uxn_opcodes_h_l654_c2_91dc_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l654_c2_91dc] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l654_c2_91dc] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l654_c2_91dc] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_cond;
     result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_return_output := result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_return_output;

     -- Submodule level 7
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l654_c2_91dc_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8040_uxn_opcodes_h_l683_l650_DUPLICATE_a750 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8040_uxn_opcodes_h_l683_l650_DUPLICATE_a750_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8040(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l654_c2_91dc_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l654_c2_91dc_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l654_c2_91dc_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l654_c2_91dc_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l654_c2_91dc_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l654_c2_91dc_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8040_uxn_opcodes_h_l683_l650_DUPLICATE_a750_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8040_uxn_opcodes_h_l683_l650_DUPLICATE_a750_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
