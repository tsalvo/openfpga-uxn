-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 52
entity and_0CLK_f62d646e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end and_0CLK_f62d646e;
architecture arch of and_0CLK_f62d646e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l947_c6_d129]
signal BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l947_c1_8811]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l947_c2_4206]
signal n8_MUX_uxn_opcodes_h_l947_c2_4206_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l947_c2_4206_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l947_c2_4206_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l947_c2_4206_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l947_c2_4206]
signal t8_MUX_uxn_opcodes_h_l947_c2_4206_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l947_c2_4206_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l947_c2_4206_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l947_c2_4206_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l947_c2_4206]
signal result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l947_c2_4206]
signal result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l947_c2_4206]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l947_c2_4206]
signal result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l947_c2_4206]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l947_c2_4206]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_return_output : unsigned(3 downto 0);

-- printf_uxn_opcodes_h_l948_c3_8e80[uxn_opcodes_h_l948_c3_8e80]
signal printf_uxn_opcodes_h_l948_c3_8e80_uxn_opcodes_h_l948_c3_8e80_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l952_c11_7d63]
signal BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l952_c7_8c18]
signal n8_MUX_uxn_opcodes_h_l952_c7_8c18_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l952_c7_8c18_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l952_c7_8c18]
signal t8_MUX_uxn_opcodes_h_l952_c7_8c18_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l952_c7_8c18_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l952_c7_8c18]
signal result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l952_c7_8c18]
signal result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l952_c7_8c18]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l952_c7_8c18]
signal result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l952_c7_8c18]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l952_c7_8c18]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l955_c11_d731]
signal BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l955_c7_72fd]
signal n8_MUX_uxn_opcodes_h_l955_c7_72fd_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l955_c7_72fd_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l955_c7_72fd]
signal t8_MUX_uxn_opcodes_h_l955_c7_72fd_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l955_c7_72fd_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l955_c7_72fd]
signal result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l955_c7_72fd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l955_c7_72fd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l955_c7_72fd]
signal result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l955_c7_72fd]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l955_c7_72fd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l959_c11_f3d1]
signal BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l959_c7_1699]
signal n8_MUX_uxn_opcodes_h_l959_c7_1699_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l959_c7_1699_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l959_c7_1699_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l959_c7_1699_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l959_c7_1699]
signal result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l959_c7_1699]
signal result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l959_c7_1699]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l959_c7_1699]
signal result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l959_c7_1699]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l959_c7_1699]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l962_c11_2af5]
signal BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l962_c7_ce3f]
signal n8_MUX_uxn_opcodes_h_l962_c7_ce3f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l962_c7_ce3f]
signal result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l962_c7_ce3f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l962_c7_ce3f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l962_c7_ce3f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l962_c7_ce3f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l962_c7_ce3f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output : unsigned(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l965_c30_5e86]
signal sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_return_output : signed(3 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l968_c21_5ad6]
signal BIN_OP_AND_uxn_opcodes_h_l968_c21_5ad6_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l968_c21_5ad6_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l968_c21_5ad6_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l970_c11_4708]
signal BIN_OP_EQ_uxn_opcodes_h_l970_c11_4708_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l970_c11_4708_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l970_c11_4708_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l970_c7_0d24]
signal result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l970_c7_0d24]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l970_c7_0d24]
signal result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_25e8( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.is_sp_shift := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129
BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_left,
BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_right,
BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_return_output);

-- n8_MUX_uxn_opcodes_h_l947_c2_4206
n8_MUX_uxn_opcodes_h_l947_c2_4206 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l947_c2_4206_cond,
n8_MUX_uxn_opcodes_h_l947_c2_4206_iftrue,
n8_MUX_uxn_opcodes_h_l947_c2_4206_iffalse,
n8_MUX_uxn_opcodes_h_l947_c2_4206_return_output);

-- t8_MUX_uxn_opcodes_h_l947_c2_4206
t8_MUX_uxn_opcodes_h_l947_c2_4206 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l947_c2_4206_cond,
t8_MUX_uxn_opcodes_h_l947_c2_4206_iftrue,
t8_MUX_uxn_opcodes_h_l947_c2_4206_iffalse,
t8_MUX_uxn_opcodes_h_l947_c2_4206_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206
result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_cond,
result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206
result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206
result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206
result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206
result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_return_output);

-- printf_uxn_opcodes_h_l948_c3_8e80_uxn_opcodes_h_l948_c3_8e80
printf_uxn_opcodes_h_l948_c3_8e80_uxn_opcodes_h_l948_c3_8e80 : entity work.printf_uxn_opcodes_h_l948_c3_8e80_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l948_c3_8e80_uxn_opcodes_h_l948_c3_8e80_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63
BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_left,
BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_right,
BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_return_output);

-- n8_MUX_uxn_opcodes_h_l952_c7_8c18
n8_MUX_uxn_opcodes_h_l952_c7_8c18 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l952_c7_8c18_cond,
n8_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue,
n8_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse,
n8_MUX_uxn_opcodes_h_l952_c7_8c18_return_output);

-- t8_MUX_uxn_opcodes_h_l952_c7_8c18
t8_MUX_uxn_opcodes_h_l952_c7_8c18 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l952_c7_8c18_cond,
t8_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue,
t8_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse,
t8_MUX_uxn_opcodes_h_l952_c7_8c18_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18
result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_cond,
result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18
result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18
result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18
result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18
result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731
BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_left,
BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_right,
BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_return_output);

-- n8_MUX_uxn_opcodes_h_l955_c7_72fd
n8_MUX_uxn_opcodes_h_l955_c7_72fd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l955_c7_72fd_cond,
n8_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue,
n8_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse,
n8_MUX_uxn_opcodes_h_l955_c7_72fd_return_output);

-- t8_MUX_uxn_opcodes_h_l955_c7_72fd
t8_MUX_uxn_opcodes_h_l955_c7_72fd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l955_c7_72fd_cond,
t8_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue,
t8_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse,
t8_MUX_uxn_opcodes_h_l955_c7_72fd_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd
result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_cond,
result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd
result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd
result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd
result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd
result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1
BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_left,
BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_right,
BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_return_output);

-- n8_MUX_uxn_opcodes_h_l959_c7_1699
n8_MUX_uxn_opcodes_h_l959_c7_1699 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l959_c7_1699_cond,
n8_MUX_uxn_opcodes_h_l959_c7_1699_iftrue,
n8_MUX_uxn_opcodes_h_l959_c7_1699_iffalse,
n8_MUX_uxn_opcodes_h_l959_c7_1699_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699
result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_cond,
result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699
result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699
result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699
result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699
result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5
BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_left,
BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_right,
BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_return_output);

-- n8_MUX_uxn_opcodes_h_l962_c7_ce3f
n8_MUX_uxn_opcodes_h_l962_c7_ce3f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l962_c7_ce3f_cond,
n8_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue,
n8_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse,
n8_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f
result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_cond,
result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f
result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f
result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f
result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f
result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output);

-- sp_relative_shift_uxn_opcodes_h_l965_c30_5e86
sp_relative_shift_uxn_opcodes_h_l965_c30_5e86 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_ins,
sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_x,
sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_y,
sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l968_c21_5ad6
BIN_OP_AND_uxn_opcodes_h_l968_c21_5ad6 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l968_c21_5ad6_left,
BIN_OP_AND_uxn_opcodes_h_l968_c21_5ad6_right,
BIN_OP_AND_uxn_opcodes_h_l968_c21_5ad6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l970_c11_4708
BIN_OP_EQ_uxn_opcodes_h_l970_c11_4708 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l970_c11_4708_left,
BIN_OP_EQ_uxn_opcodes_h_l970_c11_4708_right,
BIN_OP_EQ_uxn_opcodes_h_l970_c11_4708_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24
result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24
result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24
result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_return_output,
 n8_MUX_uxn_opcodes_h_l947_c2_4206_return_output,
 t8_MUX_uxn_opcodes_h_l947_c2_4206_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_return_output,
 n8_MUX_uxn_opcodes_h_l952_c7_8c18_return_output,
 t8_MUX_uxn_opcodes_h_l952_c7_8c18_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_return_output,
 n8_MUX_uxn_opcodes_h_l955_c7_72fd_return_output,
 t8_MUX_uxn_opcodes_h_l955_c7_72fd_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_return_output,
 n8_MUX_uxn_opcodes_h_l959_c7_1699_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_return_output,
 n8_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output,
 sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_return_output,
 BIN_OP_AND_uxn_opcodes_h_l968_c21_5ad6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l970_c11_4708_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l947_c2_4206_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l947_c2_4206_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l952_c7_8c18_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l947_c2_4206_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l947_c2_4206_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l947_c2_4206_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l947_c2_4206_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l952_c7_8c18_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l947_c2_4206_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l947_c2_4206_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l949_c3_dd41 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l948_c3_8e80_uxn_opcodes_h_l948_c3_8e80_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l955_c7_72fd_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l952_c7_8c18_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l955_c7_72fd_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l952_c7_8c18_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l953_c3_59a4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l959_c7_1699_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l955_c7_72fd_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l955_c7_72fd_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l957_c3_15f7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l959_c7_1699_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l959_c7_1699_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l959_c7_1699_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l960_c3_a1f5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l962_c7_ce3f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l967_c3_64aa : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l962_c7_ce3f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l968_c21_5ad6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l968_c21_5ad6_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l968_c21_5ad6_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l970_c11_4708_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l970_c11_4708_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l970_c11_4708_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l959_l955_l952_l947_l962_DUPLICATE_8aaf_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l959_l955_l952_l947_l962_DUPLICATE_bb98_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l959_l955_l952_l947_l970_DUPLICATE_9431_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l959_l955_l952_l947_l970_DUPLICATE_e699_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l959_l955_l952_l970_l962_DUPLICATE_3cea_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l976_l943_DUPLICATE_98be_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l970_c11_4708_right := to_unsigned(5, 3);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l953_c3_59a4 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l953_c3_59a4;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l960_c3_a1f5 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l960_c3_a1f5;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l967_c3_64aa := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l967_c3_64aa;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l957_c3_15f7 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l957_c3_15f7;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l949_c3_dd41 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l949_c3_dd41;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l947_c2_4206_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l959_c7_1699_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l970_c11_4708_left := VAR_phase;
     VAR_BIN_OP_AND_uxn_opcodes_h_l968_c21_5ad6_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_AND_uxn_opcodes_h_l968_c21_5ad6_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l947_c2_4206_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse := t8;
     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l962_c7_ce3f] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l962_c7_ce3f_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l947_c6_d129] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_left;
     BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_return_output := BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l959_l955_l952_l947_l962_DUPLICATE_bb98 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l959_l955_l952_l947_l962_DUPLICATE_bb98_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l959_l955_l952_l947_l970_DUPLICATE_e699 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l959_l955_l952_l947_l970_DUPLICATE_e699_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l955_c11_d731] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_left;
     BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_return_output := BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l968_c21_5ad6] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l968_c21_5ad6_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l968_c21_5ad6_left;
     BIN_OP_AND_uxn_opcodes_h_l968_c21_5ad6_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l968_c21_5ad6_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l968_c21_5ad6_return_output := BIN_OP_AND_uxn_opcodes_h_l968_c21_5ad6_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l959_l955_l952_l947_l962_DUPLICATE_8aaf LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l959_l955_l952_l947_l962_DUPLICATE_8aaf_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l959_c11_f3d1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_left;
     BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_return_output := BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l959_l955_l952_l947_l970_DUPLICATE_9431 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l959_l955_l952_l947_l970_DUPLICATE_9431_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l962_c11_2af5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_left;
     BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_return_output := BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l965_c30_5e86] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_ins;
     sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_x <= VAR_sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_x;
     sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_y <= VAR_sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_return_output := sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l970_c11_4708] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l970_c11_4708_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l970_c11_4708_left;
     BIN_OP_EQ_uxn_opcodes_h_l970_c11_4708_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l970_c11_4708_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l970_c11_4708_return_output := BIN_OP_EQ_uxn_opcodes_h_l970_c11_4708_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l959_l955_l952_l970_l962_DUPLICATE_3cea LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l959_l955_l952_l970_l962_DUPLICATE_3cea_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l952_c11_7d63] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_left;
     BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_return_output := BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_return_output;

     -- Submodule level 1
     VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue := VAR_BIN_OP_AND_uxn_opcodes_h_l968_c21_5ad6_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l947_c2_4206_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l947_c2_4206_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_d129_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l952_c7_8c18_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l952_c7_8c18_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_7d63_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l955_c7_72fd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l955_c7_72fd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_d731_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l959_c7_1699_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_f3d1_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l962_c7_ce3f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_2af5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l970_c11_4708_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l970_c11_4708_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l970_c11_4708_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l959_l955_l952_l947_l962_DUPLICATE_bb98_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l959_l955_l952_l947_l962_DUPLICATE_bb98_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l959_l955_l952_l947_l962_DUPLICATE_bb98_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l959_l955_l952_l947_l962_DUPLICATE_bb98_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l959_l955_l952_l947_l962_DUPLICATE_bb98_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l959_l955_l952_l970_l962_DUPLICATE_3cea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l959_l955_l952_l970_l962_DUPLICATE_3cea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l959_l955_l952_l970_l962_DUPLICATE_3cea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l959_l955_l952_l970_l962_DUPLICATE_3cea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l959_l955_l952_l970_l962_DUPLICATE_3cea_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l959_l955_l952_l947_l970_DUPLICATE_e699_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l959_l955_l952_l947_l970_DUPLICATE_e699_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l959_l955_l952_l947_l970_DUPLICATE_e699_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l959_l955_l952_l947_l970_DUPLICATE_e699_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l959_l955_l952_l947_l970_DUPLICATE_e699_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l959_l955_l952_l947_l970_DUPLICATE_9431_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l959_l955_l952_l947_l970_DUPLICATE_9431_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l959_l955_l952_l947_l970_DUPLICATE_9431_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l959_l955_l952_l947_l970_DUPLICATE_9431_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l959_l955_l952_l947_l970_DUPLICATE_9431_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l959_l955_l952_l947_l962_DUPLICATE_8aaf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l959_l955_l952_l947_l962_DUPLICATE_8aaf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l959_l955_l952_l947_l962_DUPLICATE_8aaf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l959_l955_l952_l947_l962_DUPLICATE_8aaf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l959_l955_l952_l947_l962_DUPLICATE_8aaf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l962_c7_ce3f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l965_c30_5e86_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l970_c7_0d24] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l962_c7_ce3f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l947_c1_8811] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_return_output;

     -- n8_MUX[uxn_opcodes_h_l962_c7_ce3f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l962_c7_ce3f_cond <= VAR_n8_MUX_uxn_opcodes_h_l962_c7_ce3f_cond;
     n8_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue;
     n8_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output := n8_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l962_c7_ce3f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output := result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l970_c7_0d24] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_return_output;

     -- t8_MUX[uxn_opcodes_h_l955_c7_72fd] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l955_c7_72fd_cond <= VAR_t8_MUX_uxn_opcodes_h_l955_c7_72fd_cond;
     t8_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue;
     t8_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l955_c7_72fd_return_output := t8_MUX_uxn_opcodes_h_l955_c7_72fd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l962_c7_ce3f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l970_c7_0d24] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l948_c3_8e80_uxn_opcodes_h_l948_c3_8e80_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_8811_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l959_c7_1699_iffalse := VAR_n8_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_0d24_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_0d24_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_0d24_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse := VAR_t8_MUX_uxn_opcodes_h_l955_c7_72fd_return_output;
     -- t8_MUX[uxn_opcodes_h_l952_c7_8c18] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l952_c7_8c18_cond <= VAR_t8_MUX_uxn_opcodes_h_l952_c7_8c18_cond;
     t8_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue;
     t8_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l952_c7_8c18_return_output := t8_MUX_uxn_opcodes_h_l952_c7_8c18_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l959_c7_1699] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l962_c7_ce3f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l962_c7_ce3f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output;

     -- printf_uxn_opcodes_h_l948_c3_8e80[uxn_opcodes_h_l948_c3_8e80] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l948_c3_8e80_uxn_opcodes_h_l948_c3_8e80_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l948_c3_8e80_uxn_opcodes_h_l948_c3_8e80_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_u8_value_MUX[uxn_opcodes_h_l959_c7_1699] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_cond;
     result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_return_output := result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l962_c7_ce3f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l959_c7_1699] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_return_output;

     -- n8_MUX[uxn_opcodes_h_l959_c7_1699] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l959_c7_1699_cond <= VAR_n8_MUX_uxn_opcodes_h_l959_c7_1699_cond;
     n8_MUX_uxn_opcodes_h_l959_c7_1699_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l959_c7_1699_iftrue;
     n8_MUX_uxn_opcodes_h_l959_c7_1699_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l959_c7_1699_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l959_c7_1699_return_output := n8_MUX_uxn_opcodes_h_l959_c7_1699_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse := VAR_n8_MUX_uxn_opcodes_h_l959_c7_1699_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_ce3f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_1699_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_1699_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_1699_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l947_c2_4206_iffalse := VAR_t8_MUX_uxn_opcodes_h_l952_c7_8c18_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l959_c7_1699] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l959_c7_1699] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l955_c7_72fd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_return_output;

     -- t8_MUX[uxn_opcodes_h_l947_c2_4206] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l947_c2_4206_cond <= VAR_t8_MUX_uxn_opcodes_h_l947_c2_4206_cond;
     t8_MUX_uxn_opcodes_h_l947_c2_4206_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l947_c2_4206_iftrue;
     t8_MUX_uxn_opcodes_h_l947_c2_4206_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l947_c2_4206_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l947_c2_4206_return_output := t8_MUX_uxn_opcodes_h_l947_c2_4206_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l955_c7_72fd] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_cond;
     result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_return_output := result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_return_output;

     -- n8_MUX[uxn_opcodes_h_l955_c7_72fd] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l955_c7_72fd_cond <= VAR_n8_MUX_uxn_opcodes_h_l955_c7_72fd_cond;
     n8_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue;
     n8_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l955_c7_72fd_return_output := n8_MUX_uxn_opcodes_h_l955_c7_72fd_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l955_c7_72fd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l959_c7_1699] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse := VAR_n8_MUX_uxn_opcodes_h_l955_c7_72fd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_1699_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_1699_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_1699_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_72fd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_72fd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_72fd_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l947_c2_4206_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l952_c7_8c18] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_cond;
     result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_return_output := result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_return_output;

     -- n8_MUX[uxn_opcodes_h_l952_c7_8c18] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l952_c7_8c18_cond <= VAR_n8_MUX_uxn_opcodes_h_l952_c7_8c18_cond;
     n8_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue;
     n8_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l952_c7_8c18_return_output := n8_MUX_uxn_opcodes_h_l952_c7_8c18_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l955_c7_72fd] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l952_c7_8c18] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l955_c7_72fd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l955_c7_72fd] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l952_c7_8c18] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l947_c2_4206_iffalse := VAR_n8_MUX_uxn_opcodes_h_l952_c7_8c18_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_72fd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_72fd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_72fd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8c18_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8c18_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c7_8c18_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l947_c2_4206] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l952_c7_8c18] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l952_c7_8c18] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l947_c2_4206] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l947_c2_4206] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_cond;
     result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_return_output := result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l952_c7_8c18] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_return_output;

     -- n8_MUX[uxn_opcodes_h_l947_c2_4206] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l947_c2_4206_cond <= VAR_n8_MUX_uxn_opcodes_h_l947_c2_4206_cond;
     n8_MUX_uxn_opcodes_h_l947_c2_4206_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l947_c2_4206_iftrue;
     n8_MUX_uxn_opcodes_h_l947_c2_4206_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l947_c2_4206_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l947_c2_4206_return_output := n8_MUX_uxn_opcodes_h_l947_c2_4206_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l947_c2_4206_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8c18_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8c18_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8c18_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l947_c2_4206] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l947_c2_4206] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l947_c2_4206] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l976_l943_DUPLICATE_98be LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l976_l943_DUPLICATE_98be_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_25e8(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l947_c2_4206_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_4206_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_4206_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_4206_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_4206_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_4206_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l976_l943_DUPLICATE_98be_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l976_l943_DUPLICATE_98be_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
