-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity sft_0CLK_46cced44 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sft_0CLK_46cced44;
architecture arch of sft_0CLK_46cced44 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2231_c6_179f]
signal BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2231_c2_9413]
signal t8_MUX_uxn_opcodes_h_l2231_c2_9413_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2231_c2_9413]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2231_c2_9413]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2231_c2_9413]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2231_c2_9413]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2231_c2_9413]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2231_c2_9413]
signal result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2231_c2_9413]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2231_c2_9413]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2231_c2_9413]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2231_c2_9413]
signal n8_MUX_uxn_opcodes_h_l2231_c2_9413_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2231_c2_9413]
signal tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2244_c11_fba2]
signal BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2244_c7_b7a8]
signal t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2244_c7_b7a8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2244_c7_b7a8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2244_c7_b7a8]
signal result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2244_c7_b7a8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2244_c7_b7a8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2244_c7_b7a8]
signal n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2244_c7_b7a8]
signal tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2247_c11_eee7]
signal BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2247_c7_f85b]
signal t8_MUX_uxn_opcodes_h_l2247_c7_f85b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2247_c7_f85b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2247_c7_f85b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2247_c7_f85b]
signal result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2247_c7_f85b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2247_c7_f85b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2247_c7_f85b]
signal n8_MUX_uxn_opcodes_h_l2247_c7_f85b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2247_c7_f85b]
signal tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2249_c30_e585]
signal sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2251_c11_346d]
signal BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2251_c7_9d57]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2251_c7_9d57]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2251_c7_9d57]
signal result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2251_c7_9d57]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2251_c7_9d57]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2251_c7_9d57]
signal n8_MUX_uxn_opcodes_h_l2251_c7_9d57_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2251_c7_9d57]
signal tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output : unsigned(7 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l2254_c18_9bc5]
signal BIN_OP_AND_uxn_opcodes_h_l2254_c18_9bc5_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2254_c18_9bc5_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2254_c18_9bc5_return_output : unsigned(7 downto 0);

-- BIN_OP_SR[uxn_opcodes_h_l2254_c11_f088]
signal BIN_OP_SR_uxn_opcodes_h_l2254_c11_f088_left : unsigned(7 downto 0);
signal BIN_OP_SR_uxn_opcodes_h_l2254_c11_f088_right : unsigned(7 downto 0);
signal BIN_OP_SR_uxn_opcodes_h_l2254_c11_f088_return_output : unsigned(7 downto 0);

-- CONST_SR_4[uxn_opcodes_h_l2254_c34_e6c4]
signal CONST_SR_4_uxn_opcodes_h_l2254_c34_e6c4_x : unsigned(7 downto 0);
signal CONST_SR_4_uxn_opcodes_h_l2254_c34_e6c4_return_output : unsigned(7 downto 0);

-- BIN_OP_SL[uxn_opcodes_h_l2254_c11_2006]
signal BIN_OP_SL_uxn_opcodes_h_l2254_c11_2006_left : unsigned(7 downto 0);
signal BIN_OP_SL_uxn_opcodes_h_l2254_c11_2006_right : unsigned(7 downto 0);
signal BIN_OP_SL_uxn_opcodes_h_l2254_c11_2006_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c580( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.u8_value := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_stack_index_flipped := ref_toks_8;
      base.is_pc_updated := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f
BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_left,
BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_right,
BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_return_output);

-- t8_MUX_uxn_opcodes_h_l2231_c2_9413
t8_MUX_uxn_opcodes_h_l2231_c2_9413 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2231_c2_9413_cond,
t8_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue,
t8_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse,
t8_MUX_uxn_opcodes_h_l2231_c2_9413_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413
result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413
result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413
result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413
result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413
result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_cond,
result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413
result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413
result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_return_output);

-- n8_MUX_uxn_opcodes_h_l2231_c2_9413
n8_MUX_uxn_opcodes_h_l2231_c2_9413 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2231_c2_9413_cond,
n8_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue,
n8_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse,
n8_MUX_uxn_opcodes_h_l2231_c2_9413_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2231_c2_9413
tmp8_MUX_uxn_opcodes_h_l2231_c2_9413 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_cond,
tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue,
tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse,
tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2
BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_left,
BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_right,
BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_return_output);

-- t8_MUX_uxn_opcodes_h_l2244_c7_b7a8
t8_MUX_uxn_opcodes_h_l2244_c7_b7a8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond,
t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue,
t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse,
t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8
result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8
result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond,
result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8
result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8
result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output);

-- n8_MUX_uxn_opcodes_h_l2244_c7_b7a8
n8_MUX_uxn_opcodes_h_l2244_c7_b7a8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond,
n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue,
n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse,
n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8
tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond,
tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue,
tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse,
tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7
BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_left,
BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_right,
BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_return_output);

-- t8_MUX_uxn_opcodes_h_l2247_c7_f85b
t8_MUX_uxn_opcodes_h_l2247_c7_f85b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2247_c7_f85b_cond,
t8_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue,
t8_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse,
t8_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b
result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b
result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_cond,
result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b
result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b
result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output);

-- n8_MUX_uxn_opcodes_h_l2247_c7_f85b
n8_MUX_uxn_opcodes_h_l2247_c7_f85b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2247_c7_f85b_cond,
n8_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue,
n8_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse,
n8_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b
tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_cond,
tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue,
tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse,
tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2249_c30_e585
sp_relative_shift_uxn_opcodes_h_l2249_c30_e585 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_ins,
sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_x,
sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_y,
sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d
BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_left,
BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_right,
BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57
result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57
result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_cond,
result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57
result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57
result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output);

-- n8_MUX_uxn_opcodes_h_l2251_c7_9d57
n8_MUX_uxn_opcodes_h_l2251_c7_9d57 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2251_c7_9d57_cond,
n8_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue,
n8_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse,
n8_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57
tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_cond,
tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue,
tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse,
tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l2254_c18_9bc5
BIN_OP_AND_uxn_opcodes_h_l2254_c18_9bc5 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l2254_c18_9bc5_left,
BIN_OP_AND_uxn_opcodes_h_l2254_c18_9bc5_right,
BIN_OP_AND_uxn_opcodes_h_l2254_c18_9bc5_return_output);

-- BIN_OP_SR_uxn_opcodes_h_l2254_c11_f088
BIN_OP_SR_uxn_opcodes_h_l2254_c11_f088 : entity work.BIN_OP_SR_uint8_t_uint8_t_0CLK_25d197a7 port map (
BIN_OP_SR_uxn_opcodes_h_l2254_c11_f088_left,
BIN_OP_SR_uxn_opcodes_h_l2254_c11_f088_right,
BIN_OP_SR_uxn_opcodes_h_l2254_c11_f088_return_output);

-- CONST_SR_4_uxn_opcodes_h_l2254_c34_e6c4
CONST_SR_4_uxn_opcodes_h_l2254_c34_e6c4 : entity work.CONST_SR_4_uint8_t_0CLK_de264c78 port map (
CONST_SR_4_uxn_opcodes_h_l2254_c34_e6c4_x,
CONST_SR_4_uxn_opcodes_h_l2254_c34_e6c4_return_output);

-- BIN_OP_SL_uxn_opcodes_h_l2254_c11_2006
BIN_OP_SL_uxn_opcodes_h_l2254_c11_2006 : entity work.BIN_OP_SL_uint8_t_uint8_t_0CLK_10d8c973 port map (
BIN_OP_SL_uxn_opcodes_h_l2254_c11_2006_left,
BIN_OP_SL_uxn_opcodes_h_l2254_c11_2006_right,
BIN_OP_SL_uxn_opcodes_h_l2254_c11_2006_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_return_output,
 t8_MUX_uxn_opcodes_h_l2231_c2_9413_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_return_output,
 n8_MUX_uxn_opcodes_h_l2231_c2_9413_return_output,
 tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_return_output,
 t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output,
 n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output,
 tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_return_output,
 t8_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output,
 n8_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output,
 tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output,
 sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output,
 n8_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output,
 tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output,
 BIN_OP_AND_uxn_opcodes_h_l2254_c18_9bc5_return_output,
 BIN_OP_SR_uxn_opcodes_h_l2254_c11_f088_return_output,
 CONST_SR_4_uxn_opcodes_h_l2254_c34_e6c4_return_output,
 BIN_OP_SL_uxn_opcodes_h_l2254_c11_2006_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2231_c2_9413_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2241_c3_5ea6 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2236_c3_bed4 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2231_c2_9413_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2245_c3_a1aa : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2247_c7_f85b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2247_c7_f85b_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2256_c3_7c9d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2253_c3_fcf7 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2251_c7_9d57_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2254_c11_f088_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2254_c18_9bc5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2254_c18_9bc5_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2254_c18_9bc5_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2254_c11_f088_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2254_c11_f088_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2254_c11_2006_left : unsigned(7 downto 0);
 variable VAR_CONST_SR_4_uxn_opcodes_h_l2254_c34_e6c4_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2254_c11_2006_right : unsigned(7 downto 0);
 variable VAR_CONST_SR_4_uxn_opcodes_h_l2254_c34_e6c4_x : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2254_c11_2006_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2244_l2247_l2231_l2251_DUPLICATE_3d35_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2244_l2247_l2251_DUPLICATE_dc9c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2244_l2247_l2251_DUPLICATE_a10c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2244_l2251_DUPLICATE_1518_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2247_l2251_DUPLICATE_1bf7_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l2227_l2261_DUPLICATE_c877_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_AND_uxn_opcodes_h_l2254_c18_9bc5_right := to_unsigned(15, 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_right := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_y := resize(to_signed(-1, 2), 4);
     VAR_sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2253_c3_fcf7 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2253_c3_fcf7;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2256_c3_7c9d := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2256_c3_7c9d;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2241_c3_5ea6 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2241_c3_5ea6;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2236_c3_bed4 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2236_c3_bed4;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2245_c3_a1aa := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2245_c3_a1aa;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_right := to_unsigned(3, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_left := VAR_phase;
     VAR_BIN_OP_SR_uxn_opcodes_h_l2254_c11_f088_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_AND_uxn_opcodes_h_l2254_c18_9bc5_left := t8;
     VAR_CONST_SR_4_uxn_opcodes_h_l2254_c34_e6c4_x := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse := tmp8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2231_c6_179f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2231_c2_9413] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2231_c2_9413_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2244_l2247_l2231_l2251_DUPLICATE_3d35 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2244_l2247_l2231_l2251_DUPLICATE_3d35_return_output := result.u8_value;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2231_c2_9413] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2231_c2_9413_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2247_c11_eee7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_left;
     BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_return_output := BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2231_c2_9413] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2231_c2_9413_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l2251_c11_346d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_left;
     BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_return_output := BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2244_c11_fba2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_left;
     BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_return_output := BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l2254_c18_9bc5] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l2254_c18_9bc5_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l2254_c18_9bc5_left;
     BIN_OP_AND_uxn_opcodes_h_l2254_c18_9bc5_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l2254_c18_9bc5_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l2254_c18_9bc5_return_output := BIN_OP_AND_uxn_opcodes_h_l2254_c18_9bc5_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2244_l2251_DUPLICATE_1518 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2244_l2251_DUPLICATE_1518_return_output := result.sp_relative_shift;

     -- sp_relative_shift[uxn_opcodes_h_l2249_c30_e585] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_ins;
     sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_x;
     sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_return_output := sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2244_l2247_l2251_DUPLICATE_dc9c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2244_l2247_l2251_DUPLICATE_dc9c_return_output := result.is_opc_done;

     -- CONST_SR_4[uxn_opcodes_h_l2254_c34_e6c4] LATENCY=0
     -- Inputs
     CONST_SR_4_uxn_opcodes_h_l2254_c34_e6c4_x <= VAR_CONST_SR_4_uxn_opcodes_h_l2254_c34_e6c4_x;
     -- Outputs
     VAR_CONST_SR_4_uxn_opcodes_h_l2254_c34_e6c4_return_output := CONST_SR_4_uxn_opcodes_h_l2254_c34_e6c4_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2231_c2_9413] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2231_c2_9413_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2244_l2247_l2251_DUPLICATE_a10c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2244_l2247_l2251_DUPLICATE_a10c_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2247_l2251_DUPLICATE_1bf7 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2247_l2251_DUPLICATE_1bf7_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_BIN_OP_SR_uxn_opcodes_h_l2254_c11_f088_right := VAR_BIN_OP_AND_uxn_opcodes_h_l2254_c18_9bc5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2231_c2_9413_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2231_c2_9413_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2231_c6_179f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2244_c11_fba2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2247_c7_f85b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2247_c7_f85b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2247_c11_eee7_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2251_c7_9d57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2251_c11_346d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2244_l2251_DUPLICATE_1518_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2244_l2251_DUPLICATE_1518_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2244_l2247_l2251_DUPLICATE_dc9c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2244_l2247_l2251_DUPLICATE_dc9c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2244_l2247_l2251_DUPLICATE_dc9c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2244_l2247_l2251_DUPLICATE_a10c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2244_l2247_l2251_DUPLICATE_a10c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2244_l2247_l2251_DUPLICATE_a10c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2247_l2251_DUPLICATE_1bf7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2247_l2251_DUPLICATE_1bf7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2244_l2247_l2231_l2251_DUPLICATE_3d35_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2244_l2247_l2231_l2251_DUPLICATE_3d35_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2244_l2247_l2231_l2251_DUPLICATE_3d35_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2244_l2247_l2231_l2251_DUPLICATE_3d35_return_output;
     VAR_BIN_OP_SL_uxn_opcodes_h_l2254_c11_2006_right := VAR_CONST_SR_4_uxn_opcodes_h_l2254_c34_e6c4_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2231_c2_9413_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2231_c2_9413_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2231_c2_9413_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2231_c2_9413_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2249_c30_e585_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2251_c7_9d57] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2231_c2_9413] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_return_output;

     -- BIN_OP_SR[uxn_opcodes_h_l2254_c11_f088] LATENCY=0
     -- Inputs
     BIN_OP_SR_uxn_opcodes_h_l2254_c11_f088_left <= VAR_BIN_OP_SR_uxn_opcodes_h_l2254_c11_f088_left;
     BIN_OP_SR_uxn_opcodes_h_l2254_c11_f088_right <= VAR_BIN_OP_SR_uxn_opcodes_h_l2254_c11_f088_right;
     -- Outputs
     VAR_BIN_OP_SR_uxn_opcodes_h_l2254_c11_f088_return_output := BIN_OP_SR_uxn_opcodes_h_l2254_c11_f088_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2251_c7_9d57] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output;

     -- t8_MUX[uxn_opcodes_h_l2247_c7_f85b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2247_c7_f85b_cond <= VAR_t8_MUX_uxn_opcodes_h_l2247_c7_f85b_cond;
     t8_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue;
     t8_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output := t8_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2231_c2_9413] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2251_c7_9d57] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2231_c2_9413] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2231_c2_9413] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_return_output;

     -- n8_MUX[uxn_opcodes_h_l2251_c7_9d57] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2251_c7_9d57_cond <= VAR_n8_MUX_uxn_opcodes_h_l2251_c7_9d57_cond;
     n8_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue;
     n8_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output := n8_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2251_c7_9d57] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output;

     -- Submodule level 2
     VAR_BIN_OP_SL_uxn_opcodes_h_l2254_c11_2006_left := VAR_BIN_OP_SR_uxn_opcodes_h_l2254_c11_f088_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output;
     -- t8_MUX[uxn_opcodes_h_l2244_c7_b7a8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond <= VAR_t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond;
     t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue;
     t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output := t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output;

     -- BIN_OP_SL[uxn_opcodes_h_l2254_c11_2006] LATENCY=0
     -- Inputs
     BIN_OP_SL_uxn_opcodes_h_l2254_c11_2006_left <= VAR_BIN_OP_SL_uxn_opcodes_h_l2254_c11_2006_left;
     BIN_OP_SL_uxn_opcodes_h_l2254_c11_2006_right <= VAR_BIN_OP_SL_uxn_opcodes_h_l2254_c11_2006_right;
     -- Outputs
     VAR_BIN_OP_SL_uxn_opcodes_h_l2254_c11_2006_return_output := BIN_OP_SL_uxn_opcodes_h_l2254_c11_2006_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2247_c7_f85b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2247_c7_f85b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2247_c7_f85b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output;

     -- n8_MUX[uxn_opcodes_h_l2247_c7_f85b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2247_c7_f85b_cond <= VAR_n8_MUX_uxn_opcodes_h_l2247_c7_f85b_cond;
     n8_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue;
     n8_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output := n8_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2247_c7_f85b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output;

     -- Submodule level 3
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue := VAR_BIN_OP_SL_uxn_opcodes_h_l2254_c11_2006_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue := VAR_BIN_OP_SL_uxn_opcodes_h_l2254_c11_2006_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output;
     -- t8_MUX[uxn_opcodes_h_l2231_c2_9413] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2231_c2_9413_cond <= VAR_t8_MUX_uxn_opcodes_h_l2231_c2_9413_cond;
     t8_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue;
     t8_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2231_c2_9413_return_output := t8_MUX_uxn_opcodes_h_l2231_c2_9413_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2244_c7_b7a8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2244_c7_b7a8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2251_c7_9d57] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output := result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2244_c7_b7a8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output;

     -- n8_MUX[uxn_opcodes_h_l2244_c7_b7a8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond <= VAR_n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond;
     n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue;
     n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output := n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2251_c7_9d57] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_cond;
     tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output := tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2244_c7_b7a8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2231_c2_9413_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2251_c7_9d57_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l2247_c7_f85b] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_cond;
     tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output := tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2231_c2_9413] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2231_c2_9413] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2247_c7_f85b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output := result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output;

     -- n8_MUX[uxn_opcodes_h_l2231_c2_9413] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2231_c2_9413_cond <= VAR_n8_MUX_uxn_opcodes_h_l2231_c2_9413_cond;
     n8_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue;
     n8_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2231_c2_9413_return_output := n8_MUX_uxn_opcodes_h_l2231_c2_9413_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2231_c2_9413] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2231_c2_9413] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2231_c2_9413_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2247_c7_f85b_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l2244_c7_b7a8] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond;
     tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output := tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2244_c7_b7a8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output := result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output;

     -- Submodule level 6
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2244_c7_b7a8_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2231_c2_9413] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_return_output := result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2231_c2_9413] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_cond;
     tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_return_output := tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_return_output;

     -- Submodule level 7
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l2231_c2_9413_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l2227_l2261_DUPLICATE_c877 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l2227_l2261_DUPLICATE_c877_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c580(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2231_c2_9413_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2231_c2_9413_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2231_c2_9413_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2231_c2_9413_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2231_c2_9413_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2231_c2_9413_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2231_c2_9413_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2231_c2_9413_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2231_c2_9413_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l2227_l2261_DUPLICATE_c877_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l2227_l2261_DUPLICATE_c877_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
