-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity lth_0CLK_441a128d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end lth_0CLK_441a128d;
architecture arch of lth_0CLK_441a128d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1890_c6_a527]
signal BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1890_c2_c4b9]
signal result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1890_c2_c4b9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1890_c2_c4b9]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1890_c2_c4b9]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1890_c2_c4b9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1890_c2_c4b9]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1890_c2_c4b9]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1890_c2_c4b9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1890_c2_c4b9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1890_c2_c4b9]
signal t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1890_c2_c4b9]
signal n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1903_c11_7c1b]
signal BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1903_c7_830a]
signal result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1903_c7_830a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1903_c7_830a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1903_c7_830a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1903_c7_830a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1903_c7_830a]
signal t8_MUX_uxn_opcodes_h_l1903_c7_830a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1903_c7_830a_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1903_c7_830a]
signal n8_MUX_uxn_opcodes_h_l1903_c7_830a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1903_c7_830a_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1906_c11_2c78]
signal BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1906_c7_4177]
signal result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1906_c7_4177]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1906_c7_4177]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1906_c7_4177]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1906_c7_4177]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1906_c7_4177]
signal t8_MUX_uxn_opcodes_h_l1906_c7_4177_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1906_c7_4177_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1906_c7_4177]
signal n8_MUX_uxn_opcodes_h_l1906_c7_4177_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1906_c7_4177_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1909_c11_85dd]
signal BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1909_c7_2b3b]
signal result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1909_c7_2b3b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1909_c7_2b3b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1909_c7_2b3b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1909_c7_2b3b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1909_c7_2b3b]
signal n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1911_c30_b695]
signal sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_return_output : signed(3 downto 0);

-- BIN_OP_LT[uxn_opcodes_h_l1914_c21_88f4]
signal BIN_OP_LT_uxn_opcodes_h_l1914_c21_88f4_left : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l1914_c21_88f4_right : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l1914_c21_88f4_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1914_c21_e270]
signal MUX_uxn_opcodes_h_l1914_c21_e270_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1914_c21_e270_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1914_c21_e270_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1914_c21_e270_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_243c( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : signed;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.is_vram_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_pc_updated := ref_toks_6;
      base.is_ram_write := ref_toks_7;
      base.sp_relative_shift := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527
BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_left,
BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_right,
BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9
result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond,
result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9
result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9
result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9
result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9
result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9
result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9
result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output);

-- t8_MUX_uxn_opcodes_h_l1890_c2_c4b9
t8_MUX_uxn_opcodes_h_l1890_c2_c4b9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond,
t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue,
t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse,
t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output);

-- n8_MUX_uxn_opcodes_h_l1890_c2_c4b9
n8_MUX_uxn_opcodes_h_l1890_c2_c4b9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond,
n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue,
n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse,
n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b
BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_left,
BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_right,
BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a
result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_cond,
result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a
result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a
result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a
result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_return_output);

-- t8_MUX_uxn_opcodes_h_l1903_c7_830a
t8_MUX_uxn_opcodes_h_l1903_c7_830a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1903_c7_830a_cond,
t8_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue,
t8_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse,
t8_MUX_uxn_opcodes_h_l1903_c7_830a_return_output);

-- n8_MUX_uxn_opcodes_h_l1903_c7_830a
n8_MUX_uxn_opcodes_h_l1903_c7_830a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1903_c7_830a_cond,
n8_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue,
n8_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse,
n8_MUX_uxn_opcodes_h_l1903_c7_830a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78
BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_left,
BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_right,
BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177
result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_cond,
result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177
result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177
result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177
result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_return_output);

-- t8_MUX_uxn_opcodes_h_l1906_c7_4177
t8_MUX_uxn_opcodes_h_l1906_c7_4177 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1906_c7_4177_cond,
t8_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue,
t8_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse,
t8_MUX_uxn_opcodes_h_l1906_c7_4177_return_output);

-- n8_MUX_uxn_opcodes_h_l1906_c7_4177
n8_MUX_uxn_opcodes_h_l1906_c7_4177 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1906_c7_4177_cond,
n8_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue,
n8_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse,
n8_MUX_uxn_opcodes_h_l1906_c7_4177_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd
BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd_left,
BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd_right,
BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b
result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b
result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b
result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output);

-- n8_MUX_uxn_opcodes_h_l1909_c7_2b3b
n8_MUX_uxn_opcodes_h_l1909_c7_2b3b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond,
n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue,
n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse,
n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1911_c30_b695
sp_relative_shift_uxn_opcodes_h_l1911_c30_b695 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_ins,
sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_x,
sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_y,
sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_return_output);

-- BIN_OP_LT_uxn_opcodes_h_l1914_c21_88f4
BIN_OP_LT_uxn_opcodes_h_l1914_c21_88f4 : entity work.BIN_OP_LT_uint8_t_uint8_t_0CLK_380ecc95 port map (
BIN_OP_LT_uxn_opcodes_h_l1914_c21_88f4_left,
BIN_OP_LT_uxn_opcodes_h_l1914_c21_88f4_right,
BIN_OP_LT_uxn_opcodes_h_l1914_c21_88f4_return_output);

-- MUX_uxn_opcodes_h_l1914_c21_e270
MUX_uxn_opcodes_h_l1914_c21_e270 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1914_c21_e270_cond,
MUX_uxn_opcodes_h_l1914_c21_e270_iftrue,
MUX_uxn_opcodes_h_l1914_c21_e270_iffalse,
MUX_uxn_opcodes_h_l1914_c21_e270_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output,
 t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output,
 n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_return_output,
 t8_MUX_uxn_opcodes_h_l1903_c7_830a_return_output,
 n8_MUX_uxn_opcodes_h_l1903_c7_830a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_return_output,
 t8_MUX_uxn_opcodes_h_l1906_c7_4177_return_output,
 n8_MUX_uxn_opcodes_h_l1906_c7_4177_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output,
 n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output,
 sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_return_output,
 BIN_OP_LT_uxn_opcodes_h_l1914_c21_88f4_return_output,
 MUX_uxn_opcodes_h_l1914_c21_e270_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1890_c2_c4b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1890_c2_c4b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1900_c3_8516 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1890_c2_c4b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1890_c2_c4b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1895_c3_b2a5 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1903_c7_830a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1903_c7_830a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1904_c3_c9f3 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1906_c7_4177_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1903_c7_830a_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1906_c7_4177_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1903_c7_830a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1906_c7_4177_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1906_c7_4177_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1913_c3_3101 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1914_c21_e270_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1914_c21_88f4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1914_c21_88f4_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1914_c21_88f4_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1914_c21_e270_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1914_c21_e270_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1914_c21_e270_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1906_l1890_l1909_l1903_DUPLICATE_54f1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1906_l1909_l1903_DUPLICATE_3782_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1906_l1909_l1903_DUPLICATE_3a81_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1906_l1909_l1903_DUPLICATE_f0a1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1906_l1909_DUPLICATE_82fd_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l1886_l1918_DUPLICATE_d470_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1913_c3_3101 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1913_c3_3101;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_y := resize(to_signed(-1, 2), 4);
     VAR_sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1914_c21_e270_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1895_c3_b2a5 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1895_c3_b2a5;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1904_c3_c9f3 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1904_c3_c9f3;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1900_c3_8516 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1900_c3_8516;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_right := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1914_c21_e270_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd_right := to_unsigned(3, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd_left := VAR_phase;
     VAR_BIN_OP_LT_uxn_opcodes_h_l1914_c21_88f4_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_LT_uxn_opcodes_h_l1914_c21_88f4_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse := t8;
     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1890_c2_c4b9] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1890_c2_c4b9_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1906_l1890_l1909_l1903_DUPLICATE_54f1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1906_l1890_l1909_l1903_DUPLICATE_54f1_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1909_c11_85dd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd_left;
     BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd_return_output := BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1890_c2_c4b9] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1890_c2_c4b9_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1906_l1909_l1903_DUPLICATE_3782 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1906_l1909_l1903_DUPLICATE_3782_return_output := result.is_stack_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1890_c2_c4b9] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1890_c2_c4b9_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l1903_c11_7c1b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1906_l1909_DUPLICATE_82fd LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1906_l1909_DUPLICATE_82fd_return_output := result.stack_address_sp_offset;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1890_c2_c4b9] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1890_c2_c4b9_return_output := result.is_vram_write;

     -- sp_relative_shift[uxn_opcodes_h_l1911_c30_b695] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_ins;
     sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_x;
     sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_return_output := sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_return_output;

     -- BIN_OP_LT[uxn_opcodes_h_l1914_c21_88f4] LATENCY=0
     -- Inputs
     BIN_OP_LT_uxn_opcodes_h_l1914_c21_88f4_left <= VAR_BIN_OP_LT_uxn_opcodes_h_l1914_c21_88f4_left;
     BIN_OP_LT_uxn_opcodes_h_l1914_c21_88f4_right <= VAR_BIN_OP_LT_uxn_opcodes_h_l1914_c21_88f4_right;
     -- Outputs
     VAR_BIN_OP_LT_uxn_opcodes_h_l1914_c21_88f4_return_output := BIN_OP_LT_uxn_opcodes_h_l1914_c21_88f4_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1906_l1909_l1903_DUPLICATE_f0a1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1906_l1909_l1903_DUPLICATE_f0a1_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1906_c11_2c78] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_left;
     BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_return_output := BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1906_l1909_l1903_DUPLICATE_3a81 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1906_l1909_l1903_DUPLICATE_3a81_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1890_c6_a527] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_left;
     BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_return_output := BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1890_c6_a527_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1903_c7_830a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1903_c7_830a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1903_c11_7c1b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1906_c7_4177_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1906_c7_4177_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c11_2c78_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1909_c11_85dd_return_output;
     VAR_MUX_uxn_opcodes_h_l1914_c21_e270_cond := VAR_BIN_OP_LT_uxn_opcodes_h_l1914_c21_88f4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1906_l1909_l1903_DUPLICATE_3a81_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1906_l1909_l1903_DUPLICATE_3a81_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1906_l1909_l1903_DUPLICATE_3a81_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1906_l1909_l1903_DUPLICATE_f0a1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1906_l1909_l1903_DUPLICATE_f0a1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1906_l1909_l1903_DUPLICATE_f0a1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1906_l1909_l1903_DUPLICATE_3782_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1906_l1909_l1903_DUPLICATE_3782_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1906_l1909_l1903_DUPLICATE_3782_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1906_l1909_DUPLICATE_82fd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1906_l1909_DUPLICATE_82fd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1906_l1890_l1909_l1903_DUPLICATE_54f1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1906_l1890_l1909_l1903_DUPLICATE_54f1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1906_l1890_l1909_l1903_DUPLICATE_54f1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1906_l1890_l1909_l1903_DUPLICATE_54f1_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1890_c2_c4b9_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1890_c2_c4b9_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1890_c2_c4b9_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1890_c2_c4b9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1911_c30_b695_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1909_c7_2b3b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output;

     -- MUX[uxn_opcodes_h_l1914_c21_e270] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1914_c21_e270_cond <= VAR_MUX_uxn_opcodes_h_l1914_c21_e270_cond;
     MUX_uxn_opcodes_h_l1914_c21_e270_iftrue <= VAR_MUX_uxn_opcodes_h_l1914_c21_e270_iftrue;
     MUX_uxn_opcodes_h_l1914_c21_e270_iffalse <= VAR_MUX_uxn_opcodes_h_l1914_c21_e270_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1914_c21_e270_return_output := MUX_uxn_opcodes_h_l1914_c21_e270_return_output;

     -- n8_MUX[uxn_opcodes_h_l1909_c7_2b3b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond <= VAR_n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond;
     n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue;
     n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output := n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1909_c7_2b3b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1909_c7_2b3b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output;

     -- t8_MUX[uxn_opcodes_h_l1906_c7_4177] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1906_c7_4177_cond <= VAR_t8_MUX_uxn_opcodes_h_l1906_c7_4177_cond;
     t8_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue;
     t8_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1906_c7_4177_return_output := t8_MUX_uxn_opcodes_h_l1906_c7_4177_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1890_c2_c4b9] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1890_c2_c4b9] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1909_c7_2b3b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1890_c2_c4b9] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1890_c2_c4b9] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue := VAR_MUX_uxn_opcodes_h_l1914_c21_e270_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1906_c7_4177_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1906_c7_4177] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_return_output;

     -- n8_MUX[uxn_opcodes_h_l1906_c7_4177] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1906_c7_4177_cond <= VAR_n8_MUX_uxn_opcodes_h_l1906_c7_4177_cond;
     n8_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue;
     n8_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1906_c7_4177_return_output := n8_MUX_uxn_opcodes_h_l1906_c7_4177_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1906_c7_4177] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1909_c7_2b3b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1906_c7_4177] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_return_output;

     -- t8_MUX[uxn_opcodes_h_l1903_c7_830a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1903_c7_830a_cond <= VAR_t8_MUX_uxn_opcodes_h_l1903_c7_830a_cond;
     t8_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue;
     t8_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1903_c7_830a_return_output := t8_MUX_uxn_opcodes_h_l1903_c7_830a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1906_c7_4177] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1906_c7_4177_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c7_4177_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c7_4177_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c7_4177_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c7_4177_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1909_c7_2b3b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1903_c7_830a_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1906_c7_4177] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_return_output := result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_return_output;

     -- n8_MUX[uxn_opcodes_h_l1903_c7_830a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1903_c7_830a_cond <= VAR_n8_MUX_uxn_opcodes_h_l1903_c7_830a_cond;
     n8_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue;
     n8_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1903_c7_830a_return_output := n8_MUX_uxn_opcodes_h_l1903_c7_830a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1903_c7_830a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_return_output;

     -- t8_MUX[uxn_opcodes_h_l1890_c2_c4b9] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond <= VAR_t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond;
     t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue;
     t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output := t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1903_c7_830a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1903_c7_830a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1903_c7_830a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1903_c7_830a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1903_c7_830a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1903_c7_830a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1903_c7_830a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1903_c7_830a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c7_4177_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1890_c2_c4b9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1890_c2_c4b9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1890_c2_c4b9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1903_c7_830a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_return_output := result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1890_c2_c4b9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output;

     -- n8_MUX[uxn_opcodes_h_l1890_c2_c4b9] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond <= VAR_n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond;
     n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue;
     n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output := n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1903_c7_830a_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1890_c2_c4b9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output := result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l1886_l1918_DUPLICATE_d470 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l1886_l1918_DUPLICATE_d470_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_243c(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1890_c2_c4b9_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l1886_l1918_DUPLICATE_d470_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l1886_l1918_DUPLICATE_d470_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
