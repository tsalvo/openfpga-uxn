-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 60
entity ldz2_0CLK_2ab048cc is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldz2_0CLK_2ab048cc;
architecture arch of ldz2_0CLK_2ab048cc is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8_high : unsigned(7 downto 0);
signal REG_COMB_tmp8_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1476_c6_d64d]
signal BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_return_output : unsigned(0 downto 0);

-- tmp8_high_MUX[uxn_opcodes_h_l1476_c2_6adf]
signal tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(7 downto 0);

-- tmp8_low_MUX[uxn_opcodes_h_l1476_c2_6adf]
signal tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1476_c2_6adf]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1476_c2_6adf]
signal result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1476_c2_6adf]
signal result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1476_c2_6adf]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1476_c2_6adf]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1476_c2_6adf]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1476_c2_6adf]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1476_c2_6adf]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1476_c2_6adf]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1476_c2_6adf]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1476_c2_6adf]
signal t8_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1489_c11_c786]
signal BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_return_output : unsigned(0 downto 0);

-- tmp8_high_MUX[uxn_opcodes_h_l1489_c7_f63e]
signal tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_cond : unsigned(0 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output : unsigned(7 downto 0);

-- tmp8_low_MUX[uxn_opcodes_h_l1489_c7_f63e]
signal tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_cond : unsigned(0 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1489_c7_f63e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1489_c7_f63e]
signal result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1489_c7_f63e]
signal result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1489_c7_f63e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1489_c7_f63e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1489_c7_f63e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1489_c7_f63e]
signal t8_MUX_uxn_opcodes_h_l1489_c7_f63e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1492_c11_f243]
signal BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_return_output : unsigned(0 downto 0);

-- tmp8_high_MUX[uxn_opcodes_h_l1492_c7_bca0]
signal tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_cond : unsigned(0 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output : unsigned(7 downto 0);

-- tmp8_low_MUX[uxn_opcodes_h_l1492_c7_bca0]
signal tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_cond : unsigned(0 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1492_c7_bca0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1492_c7_bca0]
signal result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1492_c7_bca0]
signal result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1492_c7_bca0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1492_c7_bca0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1492_c7_bca0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1492_c7_bca0]
signal t8_MUX_uxn_opcodes_h_l1492_c7_bca0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1494_c30_1bf6]
signal sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1497_c11_9699]
signal BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_return_output : unsigned(0 downto 0);

-- tmp8_high_MUX[uxn_opcodes_h_l1497_c7_055f]
signal tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_cond : unsigned(0 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_return_output : unsigned(7 downto 0);

-- tmp8_low_MUX[uxn_opcodes_h_l1497_c7_055f]
signal tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_cond : unsigned(0 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1497_c7_055f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1497_c7_055f]
signal result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1497_c7_055f]
signal result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1497_c7_055f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1497_c7_055f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1497_c7_055f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1499_c33_fd12]
signal BIN_OP_PLUS_uxn_opcodes_h_l1499_c33_fd12_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1499_c33_fd12_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1499_c33_fd12_return_output : unsigned(8 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1501_c11_b412]
signal BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412_return_output : unsigned(0 downto 0);

-- tmp8_high_MUX[uxn_opcodes_h_l1501_c7_780f]
signal tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_cond : unsigned(0 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_return_output : unsigned(7 downto 0);

-- tmp8_low_MUX[uxn_opcodes_h_l1501_c7_780f]
signal tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_cond : unsigned(0 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1501_c7_780f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1501_c7_780f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1501_c7_780f]
signal result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1501_c7_780f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1507_c11_e210]
signal BIN_OP_EQ_uxn_opcodes_h_l1507_c11_e210_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1507_c11_e210_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1507_c11_e210_return_output : unsigned(0 downto 0);

-- tmp8_low_MUX[uxn_opcodes_h_l1507_c7_65df]
signal tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_cond : unsigned(0 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_iftrue : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_iffalse : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1507_c7_65df]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1507_c7_65df]
signal result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1507_c7_65df]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_return_output : unsigned(0 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CAST_TO_uint16_t_uint9_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(8 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_e393( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_ram_write := ref_toks_4;
      base.is_stack_index_flipped := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_vram_write := ref_toks_8;
      base.is_pc_updated := ref_toks_9;
      base.is_opc_done := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d
BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_left,
BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_right,
BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_return_output);

-- tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf
tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_cond,
tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue,
tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse,
tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output);

-- tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf
tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_cond,
tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue,
tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse,
tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf
result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_cond,
result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf
result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_cond,
result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf
result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf
result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf
result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf
result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf
result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf
result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output);

-- t8_MUX_uxn_opcodes_h_l1476_c2_6adf
t8_MUX_uxn_opcodes_h_l1476_c2_6adf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1476_c2_6adf_cond,
t8_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue,
t8_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse,
t8_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786
BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_left,
BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_right,
BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_return_output);

-- tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e
tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_cond,
tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue,
tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse,
tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output);

-- tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e
tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_cond,
tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue,
tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse,
tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e
result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_cond,
result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e
result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_cond,
result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e
result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e
result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e
result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output);

-- t8_MUX_uxn_opcodes_h_l1489_c7_f63e
t8_MUX_uxn_opcodes_h_l1489_c7_f63e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1489_c7_f63e_cond,
t8_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue,
t8_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse,
t8_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243
BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_left,
BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_right,
BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_return_output);

-- tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0
tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_cond,
tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue,
tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse,
tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output);

-- tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0
tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_cond,
tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue,
tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse,
tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0
result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_cond,
result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0
result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_cond,
result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0
result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0
result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0
result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output);

-- t8_MUX_uxn_opcodes_h_l1492_c7_bca0
t8_MUX_uxn_opcodes_h_l1492_c7_bca0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1492_c7_bca0_cond,
t8_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue,
t8_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse,
t8_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6
sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_ins,
sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_x,
sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_y,
sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699
BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_left,
BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_right,
BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_return_output);

-- tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f
tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_cond,
tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue,
tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse,
tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_return_output);

-- tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f
tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_cond,
tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue,
tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse,
tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f
result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f
result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_cond,
result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f
result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f
result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1499_c33_fd12
BIN_OP_PLUS_uxn_opcodes_h_l1499_c33_fd12 : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1499_c33_fd12_left,
BIN_OP_PLUS_uxn_opcodes_h_l1499_c33_fd12_right,
BIN_OP_PLUS_uxn_opcodes_h_l1499_c33_fd12_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412
BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412_left,
BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412_right,
BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412_return_output);

-- tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f
tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_cond,
tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue,
tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse,
tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_return_output);

-- tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f
tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_cond,
tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue,
tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse,
tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f
result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f
result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f
result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1507_c11_e210
BIN_OP_EQ_uxn_opcodes_h_l1507_c11_e210 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1507_c11_e210_left,
BIN_OP_EQ_uxn_opcodes_h_l1507_c11_e210_right,
BIN_OP_EQ_uxn_opcodes_h_l1507_c11_e210_return_output);

-- tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df
tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_cond,
tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_iftrue,
tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_iffalse,
tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df
result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_cond,
result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df
result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8_high,
 tmp8_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_return_output,
 tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output,
 tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output,
 t8_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_return_output,
 tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output,
 tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output,
 t8_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_return_output,
 tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output,
 tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output,
 t8_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output,
 sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_return_output,
 tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_return_output,
 tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1499_c33_fd12_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412_return_output,
 tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_return_output,
 tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1507_c11_e210_return_output,
 tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1486_c3_0644 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1481_c3_8996 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1476_c2_6adf_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_cond : unsigned(0 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1490_c3_21cf : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1489_c7_f63e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_cond : unsigned(0 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1492_c7_bca0_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1495_c22_8212_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_cond : unsigned(0 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1498_c3_45ef : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1499_c33_fd12_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1499_c33_fd12_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1499_c33_fd12_return_output : unsigned(8 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1499_c22_2ed3_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_cond : unsigned(0 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1504_c3_d88e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1507_c11_e210_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1507_c11_e210_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1507_c11_e210_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1509_c3_e34d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1492_l1489_l1476_l1507_l1497_DUPLICATE_e393_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1489_l1497_l1476_DUPLICATE_1c78_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1489_l1497_l1492_l1501_DUPLICATE_1861_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1489_l1497_DUPLICATE_a1c2_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1492_l1489_l1507_l1501_l1497_DUPLICATE_92be_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1507_l1497_l1492_DUPLICATE_369d_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e393_uxn_opcodes_h_l1472_l1514_DUPLICATE_6e7d_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8_high : unsigned(7 downto 0);
variable REG_VAR_tmp8_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8_high := tmp8_high;
  REG_VAR_tmp8_low := tmp8_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1486_c3_0644 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1486_c3_0644;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1499_c33_fd12_right := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1490_c3_21cf := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1490_c3_21cf;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1481_c3_8996 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1481_c3_8996;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1498_c3_45ef := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1498_c3_45ef;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_right := to_unsigned(2, 2);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1504_c3_d88e := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1504_c3_d88e;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1507_c11_e210_right := to_unsigned(5, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1509_c3_e34d := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1509_c3_e34d;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_right := to_unsigned(3, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1507_c11_e210_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue := VAR_previous_ram_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_iftrue := VAR_previous_ram_read;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue := VAR_previous_ram_read;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1499_c33_fd12_left := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse := t8;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue := tmp8_high;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue := tmp8_high;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue := tmp8_high;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue := tmp8_high;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse := tmp8_high;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue := tmp8_low;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue := tmp8_low;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue := tmp8_low;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue := tmp8_low;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue := tmp8_low;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_iffalse := tmp8_low;
     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1489_l1497_DUPLICATE_a1c2 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1489_l1497_DUPLICATE_a1c2_return_output := result.sp_relative_shift;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1476_c2_6adf] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1476_c2_6adf_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l1489_c11_c786] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_left;
     BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_return_output := BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1499_c33_fd12] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1499_c33_fd12_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1499_c33_fd12_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1499_c33_fd12_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1499_c33_fd12_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1499_c33_fd12_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1499_c33_fd12_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1489_l1497_l1492_l1501_DUPLICATE_1861 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1489_l1497_l1492_l1501_DUPLICATE_1861_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1501_c11_b412] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412_left;
     BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412_return_output := BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1489_l1497_l1476_DUPLICATE_1c78 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1489_l1497_l1476_DUPLICATE_1c78_return_output := result.u16_value;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1507_l1497_l1492_DUPLICATE_369d LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1507_l1497_l1492_DUPLICATE_369d_return_output := result.stack_address_sp_offset;

     -- sp_relative_shift[uxn_opcodes_h_l1494_c30_1bf6] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_ins;
     sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_x;
     sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_return_output := sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1476_c2_6adf] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1476_c2_6adf_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1492_l1489_l1476_l1507_l1497_DUPLICATE_e393 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1492_l1489_l1476_l1507_l1497_DUPLICATE_e393_return_output := result.u8_value;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1495_c22_8212] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1495_c22_8212_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l1507_c11_e210] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1507_c11_e210_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1507_c11_e210_left;
     BIN_OP_EQ_uxn_opcodes_h_l1507_c11_e210_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1507_c11_e210_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1507_c11_e210_return_output := BIN_OP_EQ_uxn_opcodes_h_l1507_c11_e210_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1476_c6_d64d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1476_c2_6adf] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1476_c2_6adf_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l1492_c11_f243] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_left;
     BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_return_output := BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1476_c2_6adf] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1476_c2_6adf_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1497_c11_9699] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_left;
     BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_return_output := BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1492_l1489_l1507_l1501_l1497_DUPLICATE_92be LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1492_l1489_l1507_l1501_l1497_DUPLICATE_92be_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1476_c2_6adf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1476_c6_d64d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1489_c7_f63e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1489_c11_c786_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1492_c7_bca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1492_c11_f243_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1497_c11_9699_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1501_c11_b412_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1507_c11_e210_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1507_c11_e210_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1507_c11_e210_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1507_c11_e210_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1495_c22_8212_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1489_l1497_DUPLICATE_a1c2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1489_l1497_DUPLICATE_a1c2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1489_l1497_l1476_DUPLICATE_1c78_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1489_l1497_l1476_DUPLICATE_1c78_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1489_l1497_l1476_DUPLICATE_1c78_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1492_l1489_l1507_l1501_l1497_DUPLICATE_92be_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1492_l1489_l1507_l1501_l1497_DUPLICATE_92be_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1492_l1489_l1507_l1501_l1497_DUPLICATE_92be_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1492_l1489_l1507_l1501_l1497_DUPLICATE_92be_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1492_l1489_l1507_l1501_l1497_DUPLICATE_92be_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1489_l1497_l1492_l1501_DUPLICATE_1861_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1489_l1497_l1492_l1501_DUPLICATE_1861_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1489_l1497_l1492_l1501_DUPLICATE_1861_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1489_l1497_l1492_l1501_DUPLICATE_1861_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1507_l1497_l1492_DUPLICATE_369d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1507_l1497_l1492_DUPLICATE_369d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1507_l1497_l1492_DUPLICATE_369d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1492_l1489_l1476_l1507_l1497_DUPLICATE_e393_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1492_l1489_l1476_l1507_l1497_DUPLICATE_e393_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1492_l1489_l1476_l1507_l1497_DUPLICATE_e393_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1492_l1489_l1476_l1507_l1497_DUPLICATE_e393_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1492_l1489_l1476_l1507_l1497_DUPLICATE_e393_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1476_c2_6adf_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1476_c2_6adf_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1476_c2_6adf_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1476_c2_6adf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1494_c30_1bf6_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1507_c7_65df] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_return_output := result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_return_output;

     -- tmp8_high_MUX[uxn_opcodes_h_l1501_c7_780f] LATENCY=0
     -- Inputs
     tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_cond <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_cond;
     tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue;
     tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse;
     -- Outputs
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_return_output := tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1507_c7_65df] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_return_output;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1499_c22_2ed3] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1499_c22_2ed3_return_output := CAST_TO_uint16_t_uint9_t(
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1499_c33_fd12_return_output);

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1507_c7_65df] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_return_output;

     -- t8_MUX[uxn_opcodes_h_l1492_c7_bca0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1492_c7_bca0_cond <= VAR_t8_MUX_uxn_opcodes_h_l1492_c7_bca0_cond;
     t8_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue;
     t8_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output := t8_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1497_c7_055f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1476_c2_6adf] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output;

     -- tmp8_low_MUX[uxn_opcodes_h_l1507_c7_65df] LATENCY=0
     -- Inputs
     tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_cond <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_cond;
     tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_iftrue <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_iftrue;
     tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_iffalse <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_iffalse;
     -- Outputs
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_return_output := tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1501_c7_780f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1476_c2_6adf] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1476_c2_6adf] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1476_c2_6adf] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output;

     -- Submodule level 2
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1499_c22_2ed3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1507_c7_65df_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1501_c7_780f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1497_c7_055f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1507_c7_65df_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1507_c7_65df_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse := VAR_tmp8_high_MUX_uxn_opcodes_h_l1501_c7_780f_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse := VAR_tmp8_low_MUX_uxn_opcodes_h_l1507_c7_65df_return_output;
     -- t8_MUX[uxn_opcodes_h_l1489_c7_f63e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1489_c7_f63e_cond <= VAR_t8_MUX_uxn_opcodes_h_l1489_c7_f63e_cond;
     t8_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue;
     t8_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output := t8_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1501_c7_780f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1501_c7_780f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_return_output;

     -- tmp8_low_MUX[uxn_opcodes_h_l1501_c7_780f] LATENCY=0
     -- Inputs
     tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_cond <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_cond;
     tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue;
     tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse;
     -- Outputs
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_return_output := tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_return_output;

     -- tmp8_high_MUX[uxn_opcodes_h_l1497_c7_055f] LATENCY=0
     -- Inputs
     tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_cond <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_cond;
     tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue;
     tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse;
     -- Outputs
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_return_output := tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1501_c7_780f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1492_c7_bca0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1497_c7_055f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1497_c7_055f] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_return_output := result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1501_c7_780f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1497_c7_055f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1501_c7_780f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1497_c7_055f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1501_c7_780f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse := VAR_tmp8_high_MUX_uxn_opcodes_h_l1497_c7_055f_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse := VAR_tmp8_low_MUX_uxn_opcodes_h_l1501_c7_780f_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1497_c7_055f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1492_c7_bca0] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output := result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1497_c7_055f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_return_output;

     -- tmp8_low_MUX[uxn_opcodes_h_l1497_c7_055f] LATENCY=0
     -- Inputs
     tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_cond <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_cond;
     tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue;
     tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse;
     -- Outputs
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_return_output := tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_return_output;

     -- tmp8_high_MUX[uxn_opcodes_h_l1492_c7_bca0] LATENCY=0
     -- Inputs
     tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_cond <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_cond;
     tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue;
     tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse;
     -- Outputs
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output := tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1489_c7_f63e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1497_c7_055f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_return_output;

     -- t8_MUX[uxn_opcodes_h_l1476_c2_6adf] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1476_c2_6adf_cond <= VAR_t8_MUX_uxn_opcodes_h_l1476_c2_6adf_cond;
     t8_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue;
     t8_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output := t8_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1492_c7_bca0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1497_c7_055f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1497_c7_055f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1497_c7_055f_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse := VAR_tmp8_high_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse := VAR_tmp8_low_MUX_uxn_opcodes_h_l1497_c7_055f_return_output;
     -- tmp8_high_MUX[uxn_opcodes_h_l1489_c7_f63e] LATENCY=0
     -- Inputs
     tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_cond <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_cond;
     tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue;
     tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse;
     -- Outputs
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output := tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1489_c7_f63e] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output := result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output;

     -- tmp8_low_MUX[uxn_opcodes_h_l1492_c7_bca0] LATENCY=0
     -- Inputs
     tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_cond <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_cond;
     tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue;
     tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse;
     -- Outputs
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output := tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1492_c7_bca0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1492_c7_bca0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1476_c2_6adf] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1489_c7_f63e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1492_c7_bca0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output := result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse := VAR_tmp8_high_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse := VAR_tmp8_low_MUX_uxn_opcodes_h_l1492_c7_bca0_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1489_c7_f63e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1489_c7_f63e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output := result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1476_c2_6adf] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1489_c7_f63e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1476_c2_6adf] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output := result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output;

     -- tmp8_low_MUX[uxn_opcodes_h_l1489_c7_f63e] LATENCY=0
     -- Inputs
     tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_cond <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_cond;
     tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_iftrue;
     tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_iffalse;
     -- Outputs
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output := tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output;

     -- tmp8_high_MUX[uxn_opcodes_h_l1476_c2_6adf] LATENCY=0
     -- Inputs
     tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_cond <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_cond;
     tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue;
     tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse <= VAR_tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse;
     -- Outputs
     VAR_tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output := tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output;
     REG_VAR_tmp8_high := VAR_tmp8_high_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse := VAR_tmp8_low_MUX_uxn_opcodes_h_l1489_c7_f63e_return_output;
     -- tmp8_low_MUX[uxn_opcodes_h_l1476_c2_6adf] LATENCY=0
     -- Inputs
     tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_cond <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_cond;
     tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue;
     tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse <= VAR_tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse;
     -- Outputs
     VAR_tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output := tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1476_c2_6adf] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output := result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1476_c2_6adf] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1476_c2_6adf] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output;

     -- Submodule level 7
     REG_VAR_tmp8_low := VAR_tmp8_low_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_e393_uxn_opcodes_h_l1472_l1514_DUPLICATE_6e7d LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e393_uxn_opcodes_h_l1472_l1514_DUPLICATE_6e7d_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_e393(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1476_c2_6adf_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e393_uxn_opcodes_h_l1472_l1514_DUPLICATE_6e7d_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e393_uxn_opcodes_h_l1472_l1514_DUPLICATE_6e7d_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8_high <= REG_VAR_tmp8_high;
REG_COMB_tmp8_low <= REG_VAR_tmp8_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8_high <= REG_COMB_tmp8_high;
     tmp8_low <= REG_COMB_tmp8_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
