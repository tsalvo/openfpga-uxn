-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity gth2_0CLK_85d5529e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(15 downto 0);
 return_output : out opcode_result_t);
end gth2_0CLK_85d5529e;
architecture arch of gth2_0CLK_85d5529e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1688_c6_833c]
signal BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1688_c2_d349]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1688_c2_d349]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1688_c2_d349]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1688_c2_d349]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1688_c2_d349]
signal result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1688_c2_d349]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1688_c2_d349]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l1688_c2_d349]
signal n16_MUX_uxn_opcodes_h_l1688_c2_d349_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1688_c2_d349_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l1688_c2_d349]
signal t16_MUX_uxn_opcodes_h_l1688_c2_d349_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1688_c2_d349_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1696_c11_67b4]
signal BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1696_c7_419d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1696_c7_419d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1696_c7_419d]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1696_c7_419d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1696_c7_419d]
signal result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1696_c7_419d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1696_c7_419d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l1696_c7_419d]
signal n16_MUX_uxn_opcodes_h_l1696_c7_419d_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1696_c7_419d_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l1696_c7_419d]
signal t16_MUX_uxn_opcodes_h_l1696_c7_419d_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1696_c7_419d_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1699_c11_3f6a]
signal BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1699_c7_86d4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1699_c7_86d4]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1699_c7_86d4]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1699_c7_86d4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1699_c7_86d4]
signal result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1699_c7_86d4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1699_c7_86d4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l1699_c7_86d4]
signal n16_MUX_uxn_opcodes_h_l1699_c7_86d4_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l1699_c7_86d4]
signal t16_MUX_uxn_opcodes_h_l1699_c7_86d4_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1703_c30_e491]
signal sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1705_c11_8b98]
signal BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1705_c7_c817]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1705_c7_c817]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1705_c7_c817]
signal result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1705_c7_c817]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1705_c7_c817]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_return_output : unsigned(3 downto 0);

-- n16_MUX[uxn_opcodes_h_l1705_c7_c817]
signal n16_MUX_uxn_opcodes_h_l1705_c7_c817_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1705_c7_c817_return_output : unsigned(15 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1710_c21_2974]
signal BIN_OP_GT_uxn_opcodes_h_l1710_c21_2974_left : unsigned(15 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1710_c21_2974_right : unsigned(15 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1710_c21_2974_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1710_c21_362b]
signal MUX_uxn_opcodes_h_l1710_c21_362b_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1710_c21_362b_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1710_c21_362b_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1710_c21_362b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1712_c11_bc9f]
signal BIN_OP_EQ_uxn_opcodes_h_l1712_c11_bc9f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1712_c11_bc9f_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1712_c11_bc9f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1712_c7_ff37]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1712_c7_ff37]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_stack_operation_16bit := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_stack_write := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c
BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_left,
BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_right,
BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349
result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349
result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349
result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_cond,
result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349
result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349
result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_return_output);

-- n16_MUX_uxn_opcodes_h_l1688_c2_d349
n16_MUX_uxn_opcodes_h_l1688_c2_d349 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1688_c2_d349_cond,
n16_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue,
n16_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse,
n16_MUX_uxn_opcodes_h_l1688_c2_d349_return_output);

-- t16_MUX_uxn_opcodes_h_l1688_c2_d349
t16_MUX_uxn_opcodes_h_l1688_c2_d349 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1688_c2_d349_cond,
t16_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue,
t16_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse,
t16_MUX_uxn_opcodes_h_l1688_c2_d349_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4
BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_left,
BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_right,
BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d
result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d
result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d
result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_cond,
result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d
result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d
result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_return_output);

-- n16_MUX_uxn_opcodes_h_l1696_c7_419d
n16_MUX_uxn_opcodes_h_l1696_c7_419d : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1696_c7_419d_cond,
n16_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue,
n16_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse,
n16_MUX_uxn_opcodes_h_l1696_c7_419d_return_output);

-- t16_MUX_uxn_opcodes_h_l1696_c7_419d
t16_MUX_uxn_opcodes_h_l1696_c7_419d : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1696_c7_419d_cond,
t16_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue,
t16_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse,
t16_MUX_uxn_opcodes_h_l1696_c7_419d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a
BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_left,
BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_right,
BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4
result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4
result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4
result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_cond,
result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4
result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4
result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output);

-- n16_MUX_uxn_opcodes_h_l1699_c7_86d4
n16_MUX_uxn_opcodes_h_l1699_c7_86d4 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1699_c7_86d4_cond,
n16_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue,
n16_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse,
n16_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output);

-- t16_MUX_uxn_opcodes_h_l1699_c7_86d4
t16_MUX_uxn_opcodes_h_l1699_c7_86d4 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1699_c7_86d4_cond,
t16_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue,
t16_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse,
t16_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1703_c30_e491
sp_relative_shift_uxn_opcodes_h_l1703_c30_e491 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_ins,
sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_x,
sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_y,
sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98
BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98_left,
BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98_right,
BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817
result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817
result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817
result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_cond,
result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817
result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_return_output);

-- n16_MUX_uxn_opcodes_h_l1705_c7_c817
n16_MUX_uxn_opcodes_h_l1705_c7_c817 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1705_c7_c817_cond,
n16_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue,
n16_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse,
n16_MUX_uxn_opcodes_h_l1705_c7_c817_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1710_c21_2974
BIN_OP_GT_uxn_opcodes_h_l1710_c21_2974 : entity work.BIN_OP_GT_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1710_c21_2974_left,
BIN_OP_GT_uxn_opcodes_h_l1710_c21_2974_right,
BIN_OP_GT_uxn_opcodes_h_l1710_c21_2974_return_output);

-- MUX_uxn_opcodes_h_l1710_c21_362b
MUX_uxn_opcodes_h_l1710_c21_362b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1710_c21_362b_cond,
MUX_uxn_opcodes_h_l1710_c21_362b_iftrue,
MUX_uxn_opcodes_h_l1710_c21_362b_iffalse,
MUX_uxn_opcodes_h_l1710_c21_362b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1712_c11_bc9f
BIN_OP_EQ_uxn_opcodes_h_l1712_c11_bc9f : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1712_c11_bc9f_left,
BIN_OP_EQ_uxn_opcodes_h_l1712_c11_bc9f_right,
BIN_OP_EQ_uxn_opcodes_h_l1712_c11_bc9f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37
result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37
result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_return_output,
 n16_MUX_uxn_opcodes_h_l1688_c2_d349_return_output,
 t16_MUX_uxn_opcodes_h_l1688_c2_d349_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_return_output,
 n16_MUX_uxn_opcodes_h_l1696_c7_419d_return_output,
 t16_MUX_uxn_opcodes_h_l1696_c7_419d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output,
 n16_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output,
 t16_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output,
 sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_return_output,
 n16_MUX_uxn_opcodes_h_l1705_c7_c817_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1710_c21_2974_return_output,
 MUX_uxn_opcodes_h_l1710_c21_362b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1712_c11_bc9f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1693_c3_8ff5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1696_c7_419d_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1688_c2_d349_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1688_c2_d349_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1696_c7_419d_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1688_c2_d349_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1688_c2_d349_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1697_c3_5381 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1696_c7_419d_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1696_c7_419d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1705_c7_c817_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1699_c7_86d4_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1699_c7_86d4_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1709_c3_a9c6 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1705_c7_c817_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1710_c21_362b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1710_c21_2974_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1710_c21_2974_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1710_c21_2974_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1710_c21_362b_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1710_c21_362b_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1710_c21_362b_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1712_c11_bc9f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1712_c11_bc9f_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1712_c11_bc9f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1705_l1696_l1688_DUPLICATE_c5e5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1705_l1696_l1699_l1688_DUPLICATE_58db_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1696_l1699_l1688_DUPLICATE_fec0_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1696_l1712_l1699_l1688_DUPLICATE_2145_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1696_l1699_DUPLICATE_4409_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1705_l1696_l1712_l1699_DUPLICATE_2bd8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1705_l1699_DUPLICATE_b78a_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a_uxn_opcodes_h_l1684_l1717_DUPLICATE_4c4c_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n16 := n16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_y := resize(to_signed(-3, 3), 4);
     VAR_sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1693_c3_8ff5 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1693_c3_8ff5;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1712_c11_bc9f_right := to_unsigned(4, 3);
     VAR_MUX_uxn_opcodes_h_l1710_c21_362b_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1709_c3_a9c6 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1709_c3_a9c6;
     VAR_MUX_uxn_opcodes_h_l1710_c21_362b_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1697_c3_5381 := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1697_c3_5381;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_right := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_ins := VAR_ins;
     VAR_n16_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse := n16;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1712_c11_bc9f_left := VAR_phase;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1710_c21_2974_left := VAR_previous_stack_read;
     VAR_n16_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue := VAR_previous_stack_read;
     VAR_t16_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1710_c21_2974_right := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse := t16;
     -- BIN_OP_EQ[uxn_opcodes_h_l1688_c6_833c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1705_l1696_l1688_DUPLICATE_c5e5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1705_l1696_l1688_DUPLICATE_c5e5_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1712_c11_bc9f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1712_c11_bc9f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1712_c11_bc9f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1712_c11_bc9f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1712_c11_bc9f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1712_c11_bc9f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1712_c11_bc9f_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1703_c30_e491] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_ins;
     sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_x;
     sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_return_output := sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1696_l1699_DUPLICATE_4409 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1696_l1699_DUPLICATE_4409_return_output := result.is_stack_operation_16bit;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1696_l1699_l1688_DUPLICATE_fec0 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1696_l1699_l1688_DUPLICATE_fec0_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1696_c11_67b4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_left;
     BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_return_output := BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1705_c11_8b98] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98_left;
     BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98_return_output := BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1699_c11_3f6a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1696_l1712_l1699_l1688_DUPLICATE_2145 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1696_l1712_l1699_l1688_DUPLICATE_2145_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1705_l1699_DUPLICATE_b78a LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1705_l1699_DUPLICATE_b78a_return_output := result.stack_address_sp_offset;

     -- BIN_OP_GT[uxn_opcodes_h_l1710_c21_2974] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1710_c21_2974_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1710_c21_2974_left;
     BIN_OP_GT_uxn_opcodes_h_l1710_c21_2974_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1710_c21_2974_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1710_c21_2974_return_output := BIN_OP_GT_uxn_opcodes_h_l1710_c21_2974_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1705_l1696_l1699_l1688_DUPLICATE_58db LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1705_l1696_l1699_l1688_DUPLICATE_58db_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1705_l1696_l1712_l1699_DUPLICATE_2bd8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1705_l1696_l1712_l1699_DUPLICATE_2bd8_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_n16_MUX_uxn_opcodes_h_l1688_c2_d349_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1688_c2_d349_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1688_c6_833c_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1696_c7_419d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1696_c7_419d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1696_c11_67b4_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1699_c7_86d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1699_c7_86d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_3f6a_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1705_c7_c817_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c11_8b98_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1712_c11_bc9f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1712_c11_bc9f_return_output;
     VAR_MUX_uxn_opcodes_h_l1710_c21_362b_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1710_c21_2974_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1696_l1699_l1688_DUPLICATE_fec0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1696_l1699_l1688_DUPLICATE_fec0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1696_l1699_l1688_DUPLICATE_fec0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1705_l1696_l1712_l1699_DUPLICATE_2bd8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1705_l1696_l1712_l1699_DUPLICATE_2bd8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1705_l1696_l1712_l1699_DUPLICATE_2bd8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1705_l1696_l1712_l1699_DUPLICATE_2bd8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1705_l1696_l1688_DUPLICATE_c5e5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1705_l1696_l1688_DUPLICATE_c5e5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1705_l1696_l1688_DUPLICATE_c5e5_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1696_l1699_DUPLICATE_4409_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1696_l1699_DUPLICATE_4409_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1696_l1712_l1699_l1688_DUPLICATE_2145_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1696_l1712_l1699_l1688_DUPLICATE_2145_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1696_l1712_l1699_l1688_DUPLICATE_2145_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1696_l1712_l1699_l1688_DUPLICATE_2145_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1705_l1699_DUPLICATE_b78a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1705_l1699_DUPLICATE_b78a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1705_l1696_l1699_l1688_DUPLICATE_58db_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1705_l1696_l1699_l1688_DUPLICATE_58db_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1705_l1696_l1699_l1688_DUPLICATE_58db_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1705_l1696_l1699_l1688_DUPLICATE_58db_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1703_c30_e491_return_output;
     -- MUX[uxn_opcodes_h_l1710_c21_362b] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1710_c21_362b_cond <= VAR_MUX_uxn_opcodes_h_l1710_c21_362b_cond;
     MUX_uxn_opcodes_h_l1710_c21_362b_iftrue <= VAR_MUX_uxn_opcodes_h_l1710_c21_362b_iftrue;
     MUX_uxn_opcodes_h_l1710_c21_362b_iffalse <= VAR_MUX_uxn_opcodes_h_l1710_c21_362b_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1710_c21_362b_return_output := MUX_uxn_opcodes_h_l1710_c21_362b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1699_c7_86d4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output;

     -- t16_MUX[uxn_opcodes_h_l1699_c7_86d4] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1699_c7_86d4_cond <= VAR_t16_MUX_uxn_opcodes_h_l1699_c7_86d4_cond;
     t16_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue;
     t16_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output := t16_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output;

     -- n16_MUX[uxn_opcodes_h_l1705_c7_c817] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1705_c7_c817_cond <= VAR_n16_MUX_uxn_opcodes_h_l1705_c7_c817_cond;
     n16_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue;
     n16_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1705_c7_c817_return_output := n16_MUX_uxn_opcodes_h_l1705_c7_c817_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1699_c7_86d4] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1705_c7_c817] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1705_c7_c817] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1712_c7_ff37] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1712_c7_ff37] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue := VAR_MUX_uxn_opcodes_h_l1710_c21_362b_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1705_c7_c817_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_ff37_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1705_c7_c817_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_ff37_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c7_c817_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1705_c7_c817] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_return_output := result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_return_output;

     -- t16_MUX[uxn_opcodes_h_l1696_c7_419d] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1696_c7_419d_cond <= VAR_t16_MUX_uxn_opcodes_h_l1696_c7_419d_cond;
     t16_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue;
     t16_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1696_c7_419d_return_output := t16_MUX_uxn_opcodes_h_l1696_c7_419d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1705_c7_c817] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1696_c7_419d] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1705_c7_c817] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1699_c7_86d4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1696_c7_419d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1699_c7_86d4] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output;

     -- n16_MUX[uxn_opcodes_h_l1699_c7_86d4] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1699_c7_86d4_cond <= VAR_n16_MUX_uxn_opcodes_h_l1699_c7_86d4_cond;
     n16_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue;
     n16_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output := n16_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output;

     -- Submodule level 3
     VAR_n16_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1705_c7_c817_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1696_c7_419d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1705_c7_c817_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1696_c7_419d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1705_c7_c817_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1696_c7_419d_return_output;
     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1688_c2_d349] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_return_output;

     -- n16_MUX[uxn_opcodes_h_l1696_c7_419d] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1696_c7_419d_cond <= VAR_n16_MUX_uxn_opcodes_h_l1696_c7_419d_cond;
     n16_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue;
     n16_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1696_c7_419d_return_output := n16_MUX_uxn_opcodes_h_l1696_c7_419d_return_output;

     -- t16_MUX[uxn_opcodes_h_l1688_c2_d349] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1688_c2_d349_cond <= VAR_t16_MUX_uxn_opcodes_h_l1688_c2_d349_cond;
     t16_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue;
     t16_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1688_c2_d349_return_output := t16_MUX_uxn_opcodes_h_l1688_c2_d349_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1699_c7_86d4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1699_c7_86d4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1699_c7_86d4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output := result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1696_c7_419d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1688_c2_d349] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1696_c7_419d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_return_output;

     -- Submodule level 4
     VAR_n16_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1696_c7_419d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1696_c7_419d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1696_c7_419d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1699_c7_86d4_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l1688_c2_d349_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1688_c2_d349] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_return_output;

     -- n16_MUX[uxn_opcodes_h_l1688_c2_d349] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1688_c2_d349_cond <= VAR_n16_MUX_uxn_opcodes_h_l1688_c2_d349_cond;
     n16_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue;
     n16_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1688_c2_d349_return_output := n16_MUX_uxn_opcodes_h_l1688_c2_d349_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1696_c7_419d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1696_c7_419d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1688_c2_d349] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1696_c7_419d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_return_output := result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_return_output;

     -- Submodule level 5
     REG_VAR_n16 := VAR_n16_MUX_uxn_opcodes_h_l1688_c2_d349_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1696_c7_419d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1696_c7_419d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1696_c7_419d_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1688_c2_d349] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1688_c2_d349] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_return_output := result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1688_c2_d349] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a_uxn_opcodes_h_l1684_l1717_DUPLICATE_4c4c LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a_uxn_opcodes_h_l1684_l1717_DUPLICATE_4c4c_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1688_c2_d349_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1688_c2_d349_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1688_c2_d349_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1688_c2_d349_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1688_c2_d349_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1688_c2_d349_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1688_c2_d349_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a_uxn_opcodes_h_l1684_l1717_DUPLICATE_4c4c_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a_uxn_opcodes_h_l1684_l1717_DUPLICATE_4c4c_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n16 <= REG_VAR_n16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n16 <= REG_COMB_n16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
