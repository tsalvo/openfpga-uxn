-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity ora_0CLK_bacf6a1d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ora_0CLK_bacf6a1d;
architecture arch of ora_0CLK_bacf6a1d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l948_c6_3031]
signal BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l948_c1_e77d]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l948_c2_b990]
signal n8_MUX_uxn_opcodes_h_l948_c2_b990_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l948_c2_b990_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l948_c2_b990_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l948_c2_b990_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l948_c2_b990]
signal t8_MUX_uxn_opcodes_h_l948_c2_b990_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l948_c2_b990_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l948_c2_b990_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l948_c2_b990_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l948_c2_b990]
signal result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l948_c2_b990]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l948_c2_b990]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l948_c2_b990]
signal result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l948_c2_b990]
signal result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l948_c2_b990]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l949_c3_37d9[uxn_opcodes_h_l949_c3_37d9]
signal printf_uxn_opcodes_h_l949_c3_37d9_uxn_opcodes_h_l949_c3_37d9_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l953_c11_20c2]
signal BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l953_c7_be8d]
signal n8_MUX_uxn_opcodes_h_l953_c7_be8d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l953_c7_be8d_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l953_c7_be8d]
signal t8_MUX_uxn_opcodes_h_l953_c7_be8d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l953_c7_be8d_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l953_c7_be8d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l953_c7_be8d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l953_c7_be8d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l953_c7_be8d]
signal result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l953_c7_be8d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l953_c7_be8d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l956_c11_6d8d]
signal BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l956_c7_9580]
signal n8_MUX_uxn_opcodes_h_l956_c7_9580_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l956_c7_9580_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l956_c7_9580_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l956_c7_9580_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l956_c7_9580]
signal t8_MUX_uxn_opcodes_h_l956_c7_9580_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l956_c7_9580_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l956_c7_9580_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l956_c7_9580_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l956_c7_9580]
signal result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l956_c7_9580]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l956_c7_9580]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l956_c7_9580]
signal result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l956_c7_9580]
signal result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l956_c7_9580]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l959_c11_d4f3]
signal BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l959_c7_5d06]
signal n8_MUX_uxn_opcodes_h_l959_c7_5d06_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l959_c7_5d06_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l959_c7_5d06]
signal result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l959_c7_5d06]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l959_c7_5d06]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l959_c7_5d06]
signal result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l959_c7_5d06]
signal result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l959_c7_5d06]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l962_c30_ebf2]
signal sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_return_output : signed(3 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l965_c21_77c2]
signal BIN_OP_OR_uxn_opcodes_h_l965_c21_77c2_left : unsigned(7 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l965_c21_77c2_right : unsigned(7 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l965_c21_77c2_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l967_c11_f700]
signal BIN_OP_EQ_uxn_opcodes_h_l967_c11_f700_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l967_c11_f700_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l967_c11_f700_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l967_c7_9da7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l967_c7_9da7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l967_c7_9da7]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c551( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031
BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_left,
BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_right,
BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_return_output);

-- n8_MUX_uxn_opcodes_h_l948_c2_b990
n8_MUX_uxn_opcodes_h_l948_c2_b990 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l948_c2_b990_cond,
n8_MUX_uxn_opcodes_h_l948_c2_b990_iftrue,
n8_MUX_uxn_opcodes_h_l948_c2_b990_iffalse,
n8_MUX_uxn_opcodes_h_l948_c2_b990_return_output);

-- t8_MUX_uxn_opcodes_h_l948_c2_b990
t8_MUX_uxn_opcodes_h_l948_c2_b990 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l948_c2_b990_cond,
t8_MUX_uxn_opcodes_h_l948_c2_b990_iftrue,
t8_MUX_uxn_opcodes_h_l948_c2_b990_iffalse,
t8_MUX_uxn_opcodes_h_l948_c2_b990_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990
result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990
result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990
result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_cond,
result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990
result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990
result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_return_output);

-- printf_uxn_opcodes_h_l949_c3_37d9_uxn_opcodes_h_l949_c3_37d9
printf_uxn_opcodes_h_l949_c3_37d9_uxn_opcodes_h_l949_c3_37d9 : entity work.printf_uxn_opcodes_h_l949_c3_37d9_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l949_c3_37d9_uxn_opcodes_h_l949_c3_37d9_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2
BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_left,
BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_right,
BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_return_output);

-- n8_MUX_uxn_opcodes_h_l953_c7_be8d
n8_MUX_uxn_opcodes_h_l953_c7_be8d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l953_c7_be8d_cond,
n8_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue,
n8_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse,
n8_MUX_uxn_opcodes_h_l953_c7_be8d_return_output);

-- t8_MUX_uxn_opcodes_h_l953_c7_be8d
t8_MUX_uxn_opcodes_h_l953_c7_be8d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l953_c7_be8d_cond,
t8_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue,
t8_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse,
t8_MUX_uxn_opcodes_h_l953_c7_be8d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d
result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d
result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d
result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_cond,
result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d
result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d
result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d
BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_left,
BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_right,
BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_return_output);

-- n8_MUX_uxn_opcodes_h_l956_c7_9580
n8_MUX_uxn_opcodes_h_l956_c7_9580 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l956_c7_9580_cond,
n8_MUX_uxn_opcodes_h_l956_c7_9580_iftrue,
n8_MUX_uxn_opcodes_h_l956_c7_9580_iffalse,
n8_MUX_uxn_opcodes_h_l956_c7_9580_return_output);

-- t8_MUX_uxn_opcodes_h_l956_c7_9580
t8_MUX_uxn_opcodes_h_l956_c7_9580 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l956_c7_9580_cond,
t8_MUX_uxn_opcodes_h_l956_c7_9580_iftrue,
t8_MUX_uxn_opcodes_h_l956_c7_9580_iffalse,
t8_MUX_uxn_opcodes_h_l956_c7_9580_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580
result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580
result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_cond,
result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580
result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3
BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_left,
BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_right,
BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_return_output);

-- n8_MUX_uxn_opcodes_h_l959_c7_5d06
n8_MUX_uxn_opcodes_h_l959_c7_5d06 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l959_c7_5d06_cond,
n8_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue,
n8_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse,
n8_MUX_uxn_opcodes_h_l959_c7_5d06_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06
result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06
result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06
result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_cond,
result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06
result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06
result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_return_output);

-- sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2
sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_ins,
sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_x,
sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_y,
sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l965_c21_77c2
BIN_OP_OR_uxn_opcodes_h_l965_c21_77c2 : entity work.BIN_OP_OR_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l965_c21_77c2_left,
BIN_OP_OR_uxn_opcodes_h_l965_c21_77c2_right,
BIN_OP_OR_uxn_opcodes_h_l965_c21_77c2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l967_c11_f700
BIN_OP_EQ_uxn_opcodes_h_l967_c11_f700 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l967_c11_f700_left,
BIN_OP_EQ_uxn_opcodes_h_l967_c11_f700_right,
BIN_OP_EQ_uxn_opcodes_h_l967_c11_f700_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_return_output,
 n8_MUX_uxn_opcodes_h_l948_c2_b990_return_output,
 t8_MUX_uxn_opcodes_h_l948_c2_b990_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_return_output,
 n8_MUX_uxn_opcodes_h_l953_c7_be8d_return_output,
 t8_MUX_uxn_opcodes_h_l953_c7_be8d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_return_output,
 n8_MUX_uxn_opcodes_h_l956_c7_9580_return_output,
 t8_MUX_uxn_opcodes_h_l956_c7_9580_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_return_output,
 n8_MUX_uxn_opcodes_h_l959_c7_5d06_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_return_output,
 sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_return_output,
 BIN_OP_OR_uxn_opcodes_h_l965_c21_77c2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l967_c11_f700_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l948_c2_b990_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l948_c2_b990_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l953_c7_be8d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l948_c2_b990_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l948_c2_b990_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l948_c2_b990_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l948_c2_b990_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l953_c7_be8d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l948_c2_b990_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l948_c2_b990_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l950_c3_31bb : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l949_c3_37d9_uxn_opcodes_h_l949_c3_37d9_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l956_c7_9580_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l953_c7_be8d_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l956_c7_9580_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l953_c7_be8d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l954_c3_5805 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l956_c7_9580_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l956_c7_9580_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l959_c7_5d06_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l956_c7_9580_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l956_c7_9580_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l956_c7_9580_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l956_c7_9580_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l959_c7_5d06_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l964_c3_3745 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l965_c21_77c2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l965_c21_77c2_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l965_c21_77c2_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_f700_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_f700_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_f700_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l948_l953_l967_l956_DUPLICATE_af13_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l948_l959_l953_l956_DUPLICATE_1e9d_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l948_l959_l953_l956_DUPLICATE_c0ce_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l948_l953_l967_l956_DUPLICATE_00cf_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l959_l953_l967_l956_DUPLICATE_a7a6_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l959_l956_DUPLICATE_4be4_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l973_l944_DUPLICATE_743c_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_iftrue := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_iffalse := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l954_c3_5805 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l954_c3_5805;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_f700_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l964_c3_3745 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l964_c3_3745;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l950_c3_31bb := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l950_c3_31bb;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_right := to_unsigned(3, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l948_c2_b990_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l956_c7_9580_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_f700_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l965_c21_77c2_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l956_c7_9580_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_OR_uxn_opcodes_h_l965_c21_77c2_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l948_c2_b990_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l956_c7_9580_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l948_l953_l967_l956_DUPLICATE_af13 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l948_l953_l967_l956_DUPLICATE_af13_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l948_l959_l953_l956_DUPLICATE_c0ce LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l948_l959_l953_l956_DUPLICATE_c0ce_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l959_c11_d4f3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_left;
     BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_return_output := BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l948_l953_l967_l956_DUPLICATE_00cf LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l948_l953_l967_l956_DUPLICATE_00cf_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l956_c11_6d8d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_left;
     BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_return_output := BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l967_c11_f700] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l967_c11_f700_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_f700_left;
     BIN_OP_EQ_uxn_opcodes_h_l967_c11_f700_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_f700_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_f700_return_output := BIN_OP_EQ_uxn_opcodes_h_l967_c11_f700_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l959_l953_l967_l956_DUPLICATE_a7a6 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l959_l953_l967_l956_DUPLICATE_a7a6_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l953_c11_20c2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_left;
     BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_return_output := BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l948_c6_3031] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_left;
     BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_return_output := BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l962_c30_ebf2] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_ins;
     sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_x <= VAR_sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_x;
     sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_y <= VAR_sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_return_output := sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l948_l959_l953_l956_DUPLICATE_1e9d LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l948_l959_l953_l956_DUPLICATE_1e9d_return_output := result.sp_relative_shift;

     -- BIN_OP_OR[uxn_opcodes_h_l965_c21_77c2] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l965_c21_77c2_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l965_c21_77c2_left;
     BIN_OP_OR_uxn_opcodes_h_l965_c21_77c2_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l965_c21_77c2_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l965_c21_77c2_return_output := BIN_OP_OR_uxn_opcodes_h_l965_c21_77c2_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l959_l956_DUPLICATE_4be4 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l959_l956_DUPLICATE_4be4_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l948_c2_b990_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l948_c2_b990_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l948_c6_3031_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l953_c7_be8d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l953_c7_be8d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l953_c11_20c2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l956_c7_9580_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l956_c7_9580_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l956_c11_6d8d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l959_c7_5d06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_d4f3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_f700_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_f700_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l967_c11_f700_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l965_c21_77c2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l948_l959_l953_l956_DUPLICATE_1e9d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l948_l959_l953_l956_DUPLICATE_1e9d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l948_l959_l953_l956_DUPLICATE_1e9d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l948_l959_l953_l956_DUPLICATE_1e9d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l959_l953_l967_l956_DUPLICATE_a7a6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l959_l953_l967_l956_DUPLICATE_a7a6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l959_l953_l967_l956_DUPLICATE_a7a6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l959_l953_l967_l956_DUPLICATE_a7a6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l948_l953_l967_l956_DUPLICATE_00cf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l948_l953_l967_l956_DUPLICATE_00cf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l948_l953_l967_l956_DUPLICATE_00cf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l948_l953_l967_l956_DUPLICATE_00cf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l948_l953_l967_l956_DUPLICATE_af13_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l948_l953_l967_l956_DUPLICATE_af13_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l948_l953_l967_l956_DUPLICATE_af13_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l948_l953_l967_l956_DUPLICATE_af13_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l959_l956_DUPLICATE_4be4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l959_l956_DUPLICATE_4be4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l948_l959_l953_l956_DUPLICATE_c0ce_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l948_l959_l953_l956_DUPLICATE_c0ce_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l948_l959_l953_l956_DUPLICATE_c0ce_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l948_l959_l953_l956_DUPLICATE_c0ce_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l962_c30_ebf2_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l959_c7_5d06] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l967_c7_9da7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l959_c7_5d06] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l967_c7_9da7] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l959_c7_5d06] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_cond;
     result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_return_output := result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_return_output;

     -- t8_MUX[uxn_opcodes_h_l956_c7_9580] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l956_c7_9580_cond <= VAR_t8_MUX_uxn_opcodes_h_l956_c7_9580_cond;
     t8_MUX_uxn_opcodes_h_l956_c7_9580_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l956_c7_9580_iftrue;
     t8_MUX_uxn_opcodes_h_l956_c7_9580_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l956_c7_9580_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l956_c7_9580_return_output := t8_MUX_uxn_opcodes_h_l956_c7_9580_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l967_c7_9da7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l948_c1_e77d] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_return_output;

     -- n8_MUX[uxn_opcodes_h_l959_c7_5d06] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l959_c7_5d06_cond <= VAR_n8_MUX_uxn_opcodes_h_l959_c7_5d06_cond;
     n8_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue;
     n8_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l959_c7_5d06_return_output := n8_MUX_uxn_opcodes_h_l959_c7_5d06_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l949_c3_37d9_uxn_opcodes_h_l949_c3_37d9_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l948_c1_e77d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l956_c7_9580_iffalse := VAR_n8_MUX_uxn_opcodes_h_l959_c7_5d06_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l967_c7_9da7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l967_c7_9da7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l967_c7_9da7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_5d06_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_5d06_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_5d06_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse := VAR_t8_MUX_uxn_opcodes_h_l956_c7_9580_return_output;
     -- printf_uxn_opcodes_h_l949_c3_37d9[uxn_opcodes_h_l949_c3_37d9] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l949_c3_37d9_uxn_opcodes_h_l949_c3_37d9_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l949_c3_37d9_uxn_opcodes_h_l949_c3_37d9_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_u8_value_MUX[uxn_opcodes_h_l956_c7_9580] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_cond;
     result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_return_output := result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_return_output;

     -- t8_MUX[uxn_opcodes_h_l953_c7_be8d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l953_c7_be8d_cond <= VAR_t8_MUX_uxn_opcodes_h_l953_c7_be8d_cond;
     t8_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue;
     t8_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l953_c7_be8d_return_output := t8_MUX_uxn_opcodes_h_l953_c7_be8d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l959_c7_5d06] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l959_c7_5d06] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l959_c7_5d06] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l956_c7_9580] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_return_output;

     -- n8_MUX[uxn_opcodes_h_l956_c7_9580] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l956_c7_9580_cond <= VAR_n8_MUX_uxn_opcodes_h_l956_c7_9580_cond;
     n8_MUX_uxn_opcodes_h_l956_c7_9580_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l956_c7_9580_iftrue;
     n8_MUX_uxn_opcodes_h_l956_c7_9580_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l956_c7_9580_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l956_c7_9580_return_output := n8_MUX_uxn_opcodes_h_l956_c7_9580_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l956_c7_9580] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse := VAR_n8_MUX_uxn_opcodes_h_l956_c7_9580_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_5d06_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_5d06_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_5d06_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l956_c7_9580_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l956_c7_9580_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l956_c7_9580_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l948_c2_b990_iffalse := VAR_t8_MUX_uxn_opcodes_h_l953_c7_be8d_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l956_c7_9580] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l956_c7_9580] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l953_c7_be8d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l956_c7_9580] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l953_c7_be8d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_return_output := result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_return_output;

     -- n8_MUX[uxn_opcodes_h_l953_c7_be8d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l953_c7_be8d_cond <= VAR_n8_MUX_uxn_opcodes_h_l953_c7_be8d_cond;
     n8_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue;
     n8_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l953_c7_be8d_return_output := n8_MUX_uxn_opcodes_h_l953_c7_be8d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l953_c7_be8d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_return_output;

     -- t8_MUX[uxn_opcodes_h_l948_c2_b990] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l948_c2_b990_cond <= VAR_t8_MUX_uxn_opcodes_h_l948_c2_b990_cond;
     t8_MUX_uxn_opcodes_h_l948_c2_b990_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l948_c2_b990_iftrue;
     t8_MUX_uxn_opcodes_h_l948_c2_b990_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l948_c2_b990_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l948_c2_b990_return_output := t8_MUX_uxn_opcodes_h_l948_c2_b990_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l948_c2_b990_iffalse := VAR_n8_MUX_uxn_opcodes_h_l953_c7_be8d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l956_c7_9580_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l956_c7_9580_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l956_c7_9580_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l953_c7_be8d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l953_c7_be8d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l953_c7_be8d_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l948_c2_b990_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l953_c7_be8d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l953_c7_be8d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_return_output;

     -- n8_MUX[uxn_opcodes_h_l948_c2_b990] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l948_c2_b990_cond <= VAR_n8_MUX_uxn_opcodes_h_l948_c2_b990_cond;
     n8_MUX_uxn_opcodes_h_l948_c2_b990_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l948_c2_b990_iftrue;
     n8_MUX_uxn_opcodes_h_l948_c2_b990_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l948_c2_b990_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l948_c2_b990_return_output := n8_MUX_uxn_opcodes_h_l948_c2_b990_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l948_c2_b990] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l948_c2_b990] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_cond;
     result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_return_output := result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l953_c7_be8d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l948_c2_b990] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l948_c2_b990_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l953_c7_be8d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l953_c7_be8d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l953_c7_be8d_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l948_c2_b990] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l948_c2_b990] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l948_c2_b990] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l973_l944_DUPLICATE_743c LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l973_l944_DUPLICATE_743c_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c551(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l948_c2_b990_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l948_c2_b990_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l948_c2_b990_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l948_c2_b990_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l948_c2_b990_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l948_c2_b990_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l973_l944_DUPLICATE_743c_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l973_l944_DUPLICATE_743c_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
