-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity rot_0CLK_b288bfb7 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end rot_0CLK_b288bfb7;
architecture arch of rot_0CLK_b288bfb7 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal l8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_l8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2640_c6_97fa]
signal BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2640_c2_4da0]
signal result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2640_c2_4da0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2640_c2_4da0]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2640_c2_4da0]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2640_c2_4da0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2640_c2_4da0]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2640_c2_4da0]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2640_c2_4da0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2640_c2_4da0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2640_c2_4da0]
signal t8_MUX_uxn_opcodes_h_l2640_c2_4da0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l2640_c2_4da0]
signal l8_MUX_uxn_opcodes_h_l2640_c2_4da0_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2640_c2_4da0]
signal n8_MUX_uxn_opcodes_h_l2640_c2_4da0_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2653_c11_21f0]
signal BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2653_c7_1a43]
signal result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2653_c7_1a43]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2653_c7_1a43]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2653_c7_1a43]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2653_c7_1a43]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2653_c7_1a43]
signal t8_MUX_uxn_opcodes_h_l2653_c7_1a43_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l2653_c7_1a43]
signal l8_MUX_uxn_opcodes_h_l2653_c7_1a43_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2653_c7_1a43]
signal n8_MUX_uxn_opcodes_h_l2653_c7_1a43_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2656_c11_0def]
signal BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2656_c7_fd6d]
signal result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2656_c7_fd6d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2656_c7_fd6d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2656_c7_fd6d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2656_c7_fd6d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2656_c7_fd6d]
signal t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l2656_c7_fd6d]
signal l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2656_c7_fd6d]
signal n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2660_c11_0338]
signal BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2660_c7_7a89]
signal result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2660_c7_7a89]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2660_c7_7a89]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2660_c7_7a89]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2660_c7_7a89]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2660_c7_7a89]
signal l8_MUX_uxn_opcodes_h_l2660_c7_7a89_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2660_c7_7a89]
signal n8_MUX_uxn_opcodes_h_l2660_c7_7a89_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2662_c30_44ab]
signal sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2667_c11_0c61]
signal BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2667_c7_f698]
signal result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2667_c7_f698]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2667_c7_f698]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2667_c7_f698]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_return_output : unsigned(3 downto 0);

-- l8_MUX[uxn_opcodes_h_l2667_c7_f698]
signal l8_MUX_uxn_opcodes_h_l2667_c7_f698_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2667_c7_f698_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2673_c11_f64a]
signal BIN_OP_EQ_uxn_opcodes_h_l2673_c11_f64a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2673_c11_f64a_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2673_c11_f64a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2673_c7_bc5c]
signal result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2673_c7_bc5c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2673_c7_bc5c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_return_output : unsigned(3 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_243c( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : signed;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.is_vram_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_pc_updated := ref_toks_6;
      base.is_ram_write := ref_toks_7;
      base.sp_relative_shift := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa
BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_left,
BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_right,
BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0
result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_cond,
result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0
result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0
result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0
result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0
result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0
result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0
result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output);

-- t8_MUX_uxn_opcodes_h_l2640_c2_4da0
t8_MUX_uxn_opcodes_h_l2640_c2_4da0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2640_c2_4da0_cond,
t8_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue,
t8_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse,
t8_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output);

-- l8_MUX_uxn_opcodes_h_l2640_c2_4da0
l8_MUX_uxn_opcodes_h_l2640_c2_4da0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2640_c2_4da0_cond,
l8_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue,
l8_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse,
l8_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output);

-- n8_MUX_uxn_opcodes_h_l2640_c2_4da0
n8_MUX_uxn_opcodes_h_l2640_c2_4da0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2640_c2_4da0_cond,
n8_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue,
n8_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse,
n8_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0
BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_left,
BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_right,
BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43
result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_cond,
result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43
result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43
result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43
result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output);

-- t8_MUX_uxn_opcodes_h_l2653_c7_1a43
t8_MUX_uxn_opcodes_h_l2653_c7_1a43 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2653_c7_1a43_cond,
t8_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue,
t8_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse,
t8_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output);

-- l8_MUX_uxn_opcodes_h_l2653_c7_1a43
l8_MUX_uxn_opcodes_h_l2653_c7_1a43 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2653_c7_1a43_cond,
l8_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue,
l8_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse,
l8_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output);

-- n8_MUX_uxn_opcodes_h_l2653_c7_1a43
n8_MUX_uxn_opcodes_h_l2653_c7_1a43 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2653_c7_1a43_cond,
n8_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue,
n8_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse,
n8_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def
BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_left,
BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_right,
BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d
result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond,
result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output);

-- t8_MUX_uxn_opcodes_h_l2656_c7_fd6d
t8_MUX_uxn_opcodes_h_l2656_c7_fd6d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond,
t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue,
t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse,
t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output);

-- l8_MUX_uxn_opcodes_h_l2656_c7_fd6d
l8_MUX_uxn_opcodes_h_l2656_c7_fd6d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond,
l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue,
l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse,
l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output);

-- n8_MUX_uxn_opcodes_h_l2656_c7_fd6d
n8_MUX_uxn_opcodes_h_l2656_c7_fd6d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond,
n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue,
n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse,
n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338
BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_left,
BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_right,
BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89
result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_cond,
result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89
result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89
result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89
result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output);

-- l8_MUX_uxn_opcodes_h_l2660_c7_7a89
l8_MUX_uxn_opcodes_h_l2660_c7_7a89 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2660_c7_7a89_cond,
l8_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue,
l8_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse,
l8_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output);

-- n8_MUX_uxn_opcodes_h_l2660_c7_7a89
n8_MUX_uxn_opcodes_h_l2660_c7_7a89 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2660_c7_7a89_cond,
n8_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue,
n8_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse,
n8_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab
sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_ins,
sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_x,
sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_y,
sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61
BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61_left,
BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61_right,
BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698
result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_cond,
result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698
result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698
result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_return_output);

-- l8_MUX_uxn_opcodes_h_l2667_c7_f698
l8_MUX_uxn_opcodes_h_l2667_c7_f698 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2667_c7_f698_cond,
l8_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue,
l8_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse,
l8_MUX_uxn_opcodes_h_l2667_c7_f698_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2673_c11_f64a
BIN_OP_EQ_uxn_opcodes_h_l2673_c11_f64a : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2673_c11_f64a_left,
BIN_OP_EQ_uxn_opcodes_h_l2673_c11_f64a_right,
BIN_OP_EQ_uxn_opcodes_h_l2673_c11_f64a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 l8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output,
 t8_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output,
 l8_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output,
 n8_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output,
 t8_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output,
 l8_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output,
 n8_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output,
 t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output,
 l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output,
 n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output,
 l8_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output,
 n8_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output,
 sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_return_output,
 l8_MUX_uxn_opcodes_h_l2667_c7_f698_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2673_c11_f64a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2650_c3_fd9e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2645_c3_624d : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2640_c2_4da0_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2640_c2_4da0_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2640_c2_4da0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2654_c3_2447 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2653_c7_1a43_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2653_c7_1a43_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2653_c7_1a43_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2657_c3_5a8c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2664_c3_0a1b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2667_c7_f698_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2660_c7_7a89_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2660_c7_7a89_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2669_c3_fa07 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2670_c3_8de8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2667_c7_f698_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_f64a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_f64a_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_f64a_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2674_c3_506d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2673_c7_bc5c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2653_l2656_l2673_l2640_DUPLICATE_cfff_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2660_l2653_l2656_DUPLICATE_157b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2653_l2667_l2656_DUPLICATE_74dc_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2667_l2660_l2656_l2653_l2673_DUPLICATE_f6d3_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l2679_l2636_DUPLICATE_cc1a_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_l8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_l8 := l8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2645_c3_624d := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2645_c3_624d;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2674_c3_506d := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2674_c3_506d;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2669_c3_fa07 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2669_c3_fa07;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2650_c3_fd9e := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2650_c3_fd9e;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2657_c3_5a8c := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2657_c3_5a8c;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2654_c3_2447 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2654_c3_2447;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2670_c3_8de8 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2670_c3_8de8;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_f64a_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_right := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2664_c3_0a1b := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2664_c3_0a1b;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61_right := to_unsigned(4, 3);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_ins := VAR_ins;
     VAR_l8_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse := l8;
     VAR_n8_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_f64a_left := VAR_phase;
     VAR_l8_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse := t8;
     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2640_c2_4da0] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2640_c2_4da0_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2653_l2656_l2673_l2640_DUPLICATE_cfff LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2653_l2656_l2673_l2640_DUPLICATE_cfff_return_output := result.u8_value;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2640_c2_4da0] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2640_c2_4da0_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2660_c11_0338] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_left;
     BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_return_output := BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2667_c11_0c61] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61_left;
     BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61_return_output := BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2640_c6_97fa] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_left;
     BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_return_output := BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2662_c30_44ab] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_ins;
     sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_x;
     sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_return_output := sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2640_c2_4da0] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2640_c2_4da0_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2656_c11_0def] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_left;
     BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_return_output := BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2653_l2667_l2656_DUPLICATE_74dc LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2653_l2667_l2656_DUPLICATE_74dc_return_output := result.sp_relative_shift;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2640_c2_4da0] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2640_c2_4da0_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l2653_c11_21f0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_left;
     BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_return_output := BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2673_c11_f64a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2673_c11_f64a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_f64a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2673_c11_f64a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_f64a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_f64a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2673_c11_f64a_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2667_l2660_l2656_l2653_l2673_DUPLICATE_f6d3 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2667_l2660_l2656_l2653_l2673_DUPLICATE_f6d3_return_output := result.is_opc_done;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2673_c7_bc5c] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2673_c7_bc5c_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2660_l2653_l2656_DUPLICATE_157b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2660_l2653_l2656_DUPLICATE_157b_return_output := result.is_stack_write;

     -- Submodule level 1
     VAR_l8_MUX_uxn_opcodes_h_l2640_c2_4da0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2640_c2_4da0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2640_c2_4da0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_97fa_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2653_c7_1a43_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2653_c7_1a43_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2653_c7_1a43_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_21f0_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_0def_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2660_c7_7a89_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2660_c7_7a89_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_0338_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2667_c7_f698_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_0c61_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_f64a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_f64a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_f64a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2653_l2667_l2656_DUPLICATE_74dc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2653_l2667_l2656_DUPLICATE_74dc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2653_l2667_l2656_DUPLICATE_74dc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2667_l2660_l2656_l2653_l2673_DUPLICATE_f6d3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2667_l2660_l2656_l2653_l2673_DUPLICATE_f6d3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2667_l2660_l2656_l2653_l2673_DUPLICATE_f6d3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2667_l2660_l2656_l2653_l2673_DUPLICATE_f6d3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2667_l2660_l2656_l2653_l2673_DUPLICATE_f6d3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2660_l2653_l2656_DUPLICATE_157b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2660_l2653_l2656_DUPLICATE_157b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2660_l2653_l2656_DUPLICATE_157b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2653_l2656_l2673_l2640_DUPLICATE_cfff_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2653_l2656_l2673_l2640_DUPLICATE_cfff_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2653_l2656_l2673_l2640_DUPLICATE_cfff_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2653_l2656_l2673_l2640_DUPLICATE_cfff_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2640_c2_4da0_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2640_c2_4da0_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2640_c2_4da0_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2640_c2_4da0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2673_c7_bc5c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_44ab_return_output;
     -- result_is_vram_write_MUX[uxn_opcodes_h_l2640_c2_4da0] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2673_c7_bc5c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_return_output;

     -- n8_MUX[uxn_opcodes_h_l2660_c7_7a89] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2660_c7_7a89_cond <= VAR_n8_MUX_uxn_opcodes_h_l2660_c7_7a89_cond;
     n8_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue;
     n8_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output := n8_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2640_c2_4da0] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output;

     -- t8_MUX[uxn_opcodes_h_l2656_c7_fd6d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond <= VAR_t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond;
     t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue;
     t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output := t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2640_c2_4da0] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2673_c7_bc5c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2660_c7_7a89] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2640_c2_4da0] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2667_c7_f698] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2673_c7_bc5c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_return_output;

     -- l8_MUX[uxn_opcodes_h_l2667_c7_f698] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2667_c7_f698_cond <= VAR_l8_MUX_uxn_opcodes_h_l2667_c7_f698_cond;
     l8_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue;
     l8_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2667_c7_f698_return_output := l8_MUX_uxn_opcodes_h_l2667_c7_f698_return_output;

     -- Submodule level 2
     VAR_l8_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2667_c7_f698_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_bc5c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_f698_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_bc5c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_bc5c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2667_c7_f698] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2667_c7_f698] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_return_output := result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2667_c7_f698] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_return_output;

     -- t8_MUX[uxn_opcodes_h_l2653_c7_1a43] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2653_c7_1a43_cond <= VAR_t8_MUX_uxn_opcodes_h_l2653_c7_1a43_cond;
     t8_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue;
     t8_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output := t8_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output;

     -- n8_MUX[uxn_opcodes_h_l2656_c7_fd6d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond <= VAR_n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond;
     n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue;
     n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output := n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output;

     -- l8_MUX[uxn_opcodes_h_l2660_c7_7a89] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2660_c7_7a89_cond <= VAR_l8_MUX_uxn_opcodes_h_l2660_c7_7a89_cond;
     l8_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue;
     l8_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output := l8_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2656_c7_fd6d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2660_c7_7a89] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output;

     -- Submodule level 3
     VAR_l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_f698_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_f698_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_f698_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output;
     -- t8_MUX[uxn_opcodes_h_l2640_c2_4da0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2640_c2_4da0_cond <= VAR_t8_MUX_uxn_opcodes_h_l2640_c2_4da0_cond;
     t8_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue;
     t8_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output := t8_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output;

     -- l8_MUX[uxn_opcodes_h_l2656_c7_fd6d] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond <= VAR_l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond;
     l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue;
     l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output := l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2656_c7_fd6d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2660_c7_7a89] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output;

     -- n8_MUX[uxn_opcodes_h_l2653_c7_1a43] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2653_c7_1a43_cond <= VAR_n8_MUX_uxn_opcodes_h_l2653_c7_1a43_cond;
     n8_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue;
     n8_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output := n8_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2653_c7_1a43] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2660_c7_7a89] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2660_c7_7a89] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output := result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output;

     -- Submodule level 4
     VAR_l8_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_7a89_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2640_c2_4da0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2653_c7_1a43] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output;

     -- l8_MUX[uxn_opcodes_h_l2653_c7_1a43] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2653_c7_1a43_cond <= VAR_l8_MUX_uxn_opcodes_h_l2653_c7_1a43_cond;
     l8_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue;
     l8_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output := l8_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2656_c7_fd6d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2656_c7_fd6d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output;

     -- n8_MUX[uxn_opcodes_h_l2640_c2_4da0] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2640_c2_4da0_cond <= VAR_n8_MUX_uxn_opcodes_h_l2640_c2_4da0_cond;
     n8_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue;
     n8_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output := n8_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2656_c7_fd6d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output := result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output;

     -- Submodule level 5
     VAR_l8_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output;
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_fd6d_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2653_c7_1a43] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output := result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output;

     -- l8_MUX[uxn_opcodes_h_l2640_c2_4da0] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2640_c2_4da0_cond <= VAR_l8_MUX_uxn_opcodes_h_l2640_c2_4da0_cond;
     l8_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue;
     l8_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output := l8_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2640_c2_4da0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2653_c7_1a43] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2653_c7_1a43] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output;

     -- Submodule level 6
     REG_VAR_l8 := VAR_l8_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_1a43_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2640_c2_4da0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2640_c2_4da0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output := result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2640_c2_4da0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l2679_l2636_DUPLICATE_cc1a LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l2679_l2636_DUPLICATE_cc1a_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_243c(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_4da0_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l2679_l2636_DUPLICATE_cc1a_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l2679_l2636_DUPLICATE_cc1a_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_l8 <= REG_VAR_l8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     l8 <= REG_COMB_l8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
