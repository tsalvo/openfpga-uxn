-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 53
entity stz2_0CLK_75b4bee3 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end stz2_0CLK_75b4bee3;
architecture arch of stz2_0CLK_75b4bee3 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n16_low : unsigned(7 downto 0);
signal REG_COMB_n16_high : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1574_c6_eef0]
signal BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_return_output : unsigned(0 downto 0);

-- n16_high_MUX[uxn_opcodes_h_l1574_c2_a7d7]
signal n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1574_c2_a7d7]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1574_c2_a7d7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1574_c2_a7d7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1574_c2_a7d7]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1574_c2_a7d7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1574_c2_a7d7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1574_c2_a7d7]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1574_c2_a7d7]
signal result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1574_c2_a7d7]
signal result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(7 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1574_c2_a7d7]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(0 downto 0);

-- n16_low_MUX[uxn_opcodes_h_l1574_c2_a7d7]
signal n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1574_c2_a7d7]
signal t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1587_c11_123c]
signal BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_return_output : unsigned(0 downto 0);

-- n16_high_MUX[uxn_opcodes_h_l1587_c7_e56f]
signal n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_cond : unsigned(0 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1587_c7_e56f]
signal result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1587_c7_e56f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1587_c7_e56f]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1587_c7_e56f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1587_c7_e56f]
signal result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1587_c7_e56f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output : unsigned(3 downto 0);

-- n16_low_MUX[uxn_opcodes_h_l1587_c7_e56f]
signal n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_cond : unsigned(0 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1587_c7_e56f]
signal t8_MUX_uxn_opcodes_h_l1587_c7_e56f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1590_c11_225e]
signal BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_return_output : unsigned(0 downto 0);

-- n16_high_MUX[uxn_opcodes_h_l1590_c7_7c31]
signal n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_cond : unsigned(0 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1590_c7_7c31]
signal result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1590_c7_7c31]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1590_c7_7c31]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1590_c7_7c31]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1590_c7_7c31]
signal result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1590_c7_7c31]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output : unsigned(3 downto 0);

-- n16_low_MUX[uxn_opcodes_h_l1590_c7_7c31]
signal n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_cond : unsigned(0 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1590_c7_7c31]
signal t8_MUX_uxn_opcodes_h_l1590_c7_7c31_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1594_c11_c935]
signal BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_return_output : unsigned(0 downto 0);

-- n16_high_MUX[uxn_opcodes_h_l1594_c7_6413]
signal n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_cond : unsigned(0 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1594_c7_6413]
signal result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1594_c7_6413]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1594_c7_6413]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1594_c7_6413]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1594_c7_6413]
signal result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_return_output : unsigned(7 downto 0);

-- n16_low_MUX[uxn_opcodes_h_l1594_c7_6413]
signal n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_cond : unsigned(0 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1596_c30_09a2]
signal sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1601_c11_6ecf]
signal BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1601_c7_4b36]
signal result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1601_c7_4b36]
signal result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1601_c7_4b36]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1601_c7_4b36]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output : signed(3 downto 0);

-- n16_low_MUX[uxn_opcodes_h_l1601_c7_4b36]
signal n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_cond : unsigned(0 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output : unsigned(7 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1604_c33_8bbb]
signal BIN_OP_PLUS_uxn_opcodes_h_l1604_c33_8bbb_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1604_c33_8bbb_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1604_c33_8bbb_return_output : unsigned(8 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CAST_TO_uint16_t_uint9_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(8 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_42c1( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_ram_write := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_index_flipped := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.u16_value := ref_toks_8;
      base.u8_value := ref_toks_9;
      base.is_vram_write := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0
BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_left,
BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_right,
BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_return_output);

-- n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7
n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond,
n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue,
n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse,
n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7
result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7
result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7
result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7
result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7
result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7
result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond,
result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7
result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond,
result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7
result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output);

-- n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7
n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond,
n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue,
n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse,
n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output);

-- t8_MUX_uxn_opcodes_h_l1574_c2_a7d7
t8_MUX_uxn_opcodes_h_l1574_c2_a7d7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond,
t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue,
t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse,
t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c
BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_left,
BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_right,
BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_return_output);

-- n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f
n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_cond,
n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue,
n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse,
n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f
result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_cond,
result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f
result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f
result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f
result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output);

-- n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f
n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_cond,
n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue,
n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse,
n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output);

-- t8_MUX_uxn_opcodes_h_l1587_c7_e56f
t8_MUX_uxn_opcodes_h_l1587_c7_e56f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1587_c7_e56f_cond,
t8_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue,
t8_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse,
t8_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e
BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_left,
BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_right,
BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_return_output);

-- n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31
n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_cond,
n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue,
n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse,
n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31
result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_cond,
result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31
result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31
result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31
result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31
result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_cond,
result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output);

-- n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31
n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_cond,
n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue,
n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse,
n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output);

-- t8_MUX_uxn_opcodes_h_l1590_c7_7c31
t8_MUX_uxn_opcodes_h_l1590_c7_7c31 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1590_c7_7c31_cond,
t8_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue,
t8_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse,
t8_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935
BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_left,
BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_right,
BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_return_output);

-- n16_high_MUX_uxn_opcodes_h_l1594_c7_6413
n16_high_MUX_uxn_opcodes_h_l1594_c7_6413 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_cond,
n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue,
n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse,
n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413
result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_cond,
result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413
result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413
result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413
result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413
result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_cond,
result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_return_output);

-- n16_low_MUX_uxn_opcodes_h_l1594_c7_6413
n16_low_MUX_uxn_opcodes_h_l1594_c7_6413 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_cond,
n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue,
n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse,
n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2
sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_ins,
sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_x,
sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_y,
sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf
BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf_left,
BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf_right,
BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36
result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_cond,
result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36
result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_cond,
result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36
result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36
result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output);

-- n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36
n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_cond,
n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue,
n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse,
n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1604_c33_8bbb
BIN_OP_PLUS_uxn_opcodes_h_l1604_c33_8bbb : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1604_c33_8bbb_left,
BIN_OP_PLUS_uxn_opcodes_h_l1604_c33_8bbb_right,
BIN_OP_PLUS_uxn_opcodes_h_l1604_c33_8bbb_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n16_low,
 n16_high,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_return_output,
 n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output,
 n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output,
 t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_return_output,
 n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output,
 n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output,
 t8_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_return_output,
 n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output,
 n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output,
 t8_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_return_output,
 n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_return_output,
 n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_return_output,
 sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output,
 n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1604_c33_8bbb_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_return_output : unsigned(0 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1579_c3_d154 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1584_c3_0a39 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_return_output : unsigned(0 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1588_c3_6f07 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_cond : unsigned(0 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1587_c7_e56f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_return_output : unsigned(0 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_return_output : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1592_c3_8413 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1590_c7_7c31_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_cond : unsigned(0 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_return_output : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1590_c7_7c31_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_return_output : unsigned(0 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_cond : unsigned(0 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1598_c22_de93_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1603_c3_d7fa : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_cond : unsigned(0 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1604_c33_8bbb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1604_c33_8bbb_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1604_c33_8bbb_return_output : unsigned(8 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1604_c22_ea21_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1587_l1601_l1590_l1574_DUPLICATE_bc6c_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1587_l1601_l1590_l1574_DUPLICATE_f1ff_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1587_l1594_l1590_l1601_DUPLICATE_5e2f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1587_l1594_l1590_DUPLICATE_a009_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1587_l1590_l1601_DUPLICATE_4b22_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_42c1_uxn_opcodes_h_l1609_l1569_DUPLICATE_287e_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n16_low : unsigned(7 downto 0);
variable REG_VAR_n16_high : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n16_low := n16_low;
  REG_VAR_n16_high := n16_high;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf_right := to_unsigned(4, 3);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1579_c3_d154 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1579_c3_d154;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1592_c3_8413 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1592_c3_8413;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_right := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1604_c33_8bbb_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_y := resize(to_signed(-3, 3), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_right := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1588_c3_6f07 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1588_c3_6f07;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1603_c3_d7fa := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1603_c3_d7fa;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1584_c3_0a39 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1584_c3_0a39;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_ins := VAR_ins;
     VAR_n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue := n16_high;
     VAR_n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue := n16_high;
     VAR_n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue := n16_high;
     VAR_n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse := n16_high;
     VAR_n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue := n16_low;
     VAR_n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue := n16_low;
     VAR_n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue := n16_low;
     VAR_n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue := n16_low;
     VAR_n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse := n16_low;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf_left := VAR_phase;
     VAR_n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue := VAR_previous_stack_read;
     VAR_n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1604_c33_8bbb_left := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse := t8;
     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1587_l1601_l1590_l1574_DUPLICATE_f1ff LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1587_l1601_l1590_l1574_DUPLICATE_f1ff_return_output := result.u8_value;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1574_c2_a7d7] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1574_c2_a7d7_return_output := result.is_vram_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1587_l1590_l1601_DUPLICATE_4b22 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1587_l1590_l1601_DUPLICATE_4b22_return_output := result.sp_relative_shift;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1598_c22_de93] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1598_c22_de93_return_output := CAST_TO_uint16_t_uint8_t(
     t8);

     -- BIN_OP_EQ[uxn_opcodes_h_l1601_c11_6ecf] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf_left;
     BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf_return_output := BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1590_c7_7c31] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1590_c7_7c31_return_output := result.stack_address_sp_offset;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1574_c2_a7d7] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1574_c2_a7d7_return_output := result.is_pc_updated;

     -- result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d[uxn_opcodes_h_l1574_c2_a7d7] LATENCY=0
     VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1574_c2_a7d7_return_output := result.is_stack_write;

     -- sp_relative_shift[uxn_opcodes_h_l1596_c30_09a2] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_ins;
     sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_x;
     sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_return_output := sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1587_l1594_l1590_DUPLICATE_a009 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1587_l1594_l1590_DUPLICATE_a009_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1587_c11_123c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1604_c33_8bbb] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1604_c33_8bbb_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1604_c33_8bbb_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1604_c33_8bbb_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1604_c33_8bbb_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1604_c33_8bbb_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1604_c33_8bbb_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1587_l1594_l1590_l1601_DUPLICATE_5e2f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1587_l1594_l1590_l1601_DUPLICATE_5e2f_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1594_c11_c935] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_left;
     BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_return_output := BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1574_c6_eef0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_left;
     BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_return_output := BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1590_c11_225e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1587_l1601_l1590_l1574_DUPLICATE_bc6c LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1587_l1601_l1590_l1574_DUPLICATE_bc6c_return_output := result.u16_value;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1574_c2_a7d7] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1574_c2_a7d7_return_output := result.is_stack_index_flipped;

     -- Submodule level 1
     VAR_n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1574_c6_eef0_return_output;
     VAR_n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1587_c7_e56f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1587_c11_123c_return_output;
     VAR_n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1590_c7_7c31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1590_c11_225e_return_output;
     VAR_n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1594_c11_c935_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1601_c11_6ecf_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1598_c22_de93_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1587_l1590_l1601_DUPLICATE_4b22_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1587_l1590_l1601_DUPLICATE_4b22_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1587_l1590_l1601_DUPLICATE_4b22_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1587_l1601_l1590_l1574_DUPLICATE_bc6c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1587_l1601_l1590_l1574_DUPLICATE_bc6c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1587_l1601_l1590_l1574_DUPLICATE_bc6c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1587_l1601_l1590_l1574_DUPLICATE_bc6c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1587_l1594_l1590_l1601_DUPLICATE_5e2f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1587_l1594_l1590_l1601_DUPLICATE_5e2f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1587_l1594_l1590_l1601_DUPLICATE_5e2f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1587_l1594_l1590_l1601_DUPLICATE_5e2f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1587_l1594_l1590_DUPLICATE_a009_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1587_l1594_l1590_DUPLICATE_a009_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1587_l1594_l1590_DUPLICATE_a009_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1587_l1601_l1590_l1574_DUPLICATE_f1ff_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1587_l1601_l1590_l1574_DUPLICATE_f1ff_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1587_l1601_l1590_l1574_DUPLICATE_f1ff_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1587_l1601_l1590_l1574_DUPLICATE_f1ff_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1574_c2_a7d7_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1574_c2_a7d7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse := VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1574_c2_a7d7_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1574_c2_a7d7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1590_c7_7c31_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1596_c30_09a2_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1601_c7_4b36] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output;

     -- n16_high_MUX[uxn_opcodes_h_l1594_c7_6413] LATENCY=0
     -- Inputs
     n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_cond <= VAR_n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_cond;
     n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue <= VAR_n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue;
     n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse <= VAR_n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse;
     -- Outputs
     VAR_n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_return_output := n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_return_output;

     -- n16_low_MUX[uxn_opcodes_h_l1601_c7_4b36] LATENCY=0
     -- Inputs
     n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_cond <= VAR_n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_cond;
     n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue <= VAR_n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue;
     n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse <= VAR_n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse;
     -- Outputs
     VAR_n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output := n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1594_c7_6413] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1574_c2_a7d7] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1574_c2_a7d7] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1590_c7_7c31] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1574_c2_a7d7] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1601_c7_4b36] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output := result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1574_c2_a7d7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output;

     -- t8_MUX[uxn_opcodes_h_l1590_c7_7c31] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1590_c7_7c31_cond <= VAR_t8_MUX_uxn_opcodes_h_l1590_c7_7c31_cond;
     t8_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue;
     t8_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output := t8_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1604_c22_ea21] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1604_c22_ea21_return_output := CAST_TO_uint16_t_uint9_t(
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1604_c33_8bbb_return_output);

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1601_c7_4b36] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output;

     -- Submodule level 2
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1604_c22_ea21_return_output;
     VAR_n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse := VAR_n16_high_MUX_uxn_opcodes_h_l1594_c7_6413_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse := VAR_n16_low_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1594_c7_6413_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output;
     -- result_is_ram_write_MUX[uxn_opcodes_h_l1590_c7_7c31] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output;

     -- t8_MUX[uxn_opcodes_h_l1587_c7_e56f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1587_c7_e56f_cond <= VAR_t8_MUX_uxn_opcodes_h_l1587_c7_e56f_cond;
     t8_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue;
     t8_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output := t8_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output;

     -- n16_high_MUX[uxn_opcodes_h_l1590_c7_7c31] LATENCY=0
     -- Inputs
     n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_cond <= VAR_n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_cond;
     n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue <= VAR_n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue;
     n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse <= VAR_n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse;
     -- Outputs
     VAR_n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output := n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1594_c7_6413] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1594_c7_6413] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1587_c7_e56f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1601_c7_4b36] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output := result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1594_c7_6413] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_return_output := result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_return_output;

     -- n16_low_MUX[uxn_opcodes_h_l1594_c7_6413] LATENCY=0
     -- Inputs
     n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_cond <= VAR_n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_cond;
     n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue <= VAR_n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue;
     n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse <= VAR_n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse;
     -- Outputs
     VAR_n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_return_output := n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_return_output;

     -- Submodule level 3
     VAR_n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse := VAR_n16_high_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse := VAR_n16_low_MUX_uxn_opcodes_h_l1594_c7_6413_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1594_c7_6413_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1594_c7_6413_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1601_c7_4b36_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1594_c7_6413_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1590_c7_7c31] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output := result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1594_c7_6413] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_return_output := result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1590_c7_7c31] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output;

     -- n16_high_MUX[uxn_opcodes_h_l1587_c7_e56f] LATENCY=0
     -- Inputs
     n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_cond <= VAR_n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_cond;
     n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue <= VAR_n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue;
     n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse <= VAR_n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse;
     -- Outputs
     VAR_n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output := n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output;

     -- t8_MUX[uxn_opcodes_h_l1574_c2_a7d7] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond <= VAR_t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond;
     t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue;
     t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output := t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output;

     -- n16_low_MUX[uxn_opcodes_h_l1590_c7_7c31] LATENCY=0
     -- Inputs
     n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_cond <= VAR_n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_cond;
     n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue <= VAR_n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue;
     n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse <= VAR_n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse;
     -- Outputs
     VAR_n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output := n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1587_c7_e56f] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1590_c7_7c31] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1574_c2_a7d7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output;

     -- Submodule level 4
     VAR_n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse := VAR_n16_high_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse := VAR_n16_low_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1594_c7_6413_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output;
     -- n16_high_MUX[uxn_opcodes_h_l1574_c2_a7d7] LATENCY=0
     -- Inputs
     n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond <= VAR_n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond;
     n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue <= VAR_n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue;
     n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse <= VAR_n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse;
     -- Outputs
     VAR_n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output := n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1587_c7_e56f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1587_c7_e56f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1587_c7_e56f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1574_c2_a7d7] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1590_c7_7c31] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output := result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output;

     -- n16_low_MUX[uxn_opcodes_h_l1587_c7_e56f] LATENCY=0
     -- Inputs
     n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_cond <= VAR_n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_cond;
     n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue <= VAR_n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue;
     n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse <= VAR_n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse;
     -- Outputs
     VAR_n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output := n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output;

     -- Submodule level 5
     REG_VAR_n16_high := VAR_n16_high_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse := VAR_n16_low_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1590_c7_7c31_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output;
     -- n16_low_MUX[uxn_opcodes_h_l1574_c2_a7d7] LATENCY=0
     -- Inputs
     n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond <= VAR_n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond;
     n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue <= VAR_n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue;
     n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse <= VAR_n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse;
     -- Outputs
     VAR_n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output := n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1574_c2_a7d7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1574_c2_a7d7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output := result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1574_c2_a7d7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1587_c7_e56f] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output := result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output;

     -- Submodule level 6
     REG_VAR_n16_low := VAR_n16_low_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1587_c7_e56f_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l1574_c2_a7d7] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output := result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_42c1_uxn_opcodes_h_l1609_l1569_DUPLICATE_287e LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_42c1_uxn_opcodes_h_l1609_l1569_DUPLICATE_287e_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_42c1(
     result,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1574_c2_a7d7_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_42c1_uxn_opcodes_h_l1609_l1569_DUPLICATE_287e_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_42c1_uxn_opcodes_h_l1609_l1569_DUPLICATE_287e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n16_low <= REG_VAR_n16_low;
REG_COMB_n16_high <= REG_VAR_n16_high;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n16_low <= REG_COMB_n16_low;
     n16_high <= REG_COMB_n16_high;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
