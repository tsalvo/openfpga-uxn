-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity neq_0CLK_85d5529e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end neq_0CLK_85d5529e;
architecture arch of neq_0CLK_85d5529e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1188_c6_7c4d]
signal BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1188_c1_afa1]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1188_c2_5b1f]
signal t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1188_c2_5b1f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1188_c2_5b1f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1188_c2_5b1f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1188_c2_5b1f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1188_c2_5b1f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1188_c2_5b1f]
signal result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1188_c2_5b1f]
signal n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1189_c3_f7be[uxn_opcodes_h_l1189_c3_f7be]
signal printf_uxn_opcodes_h_l1189_c3_f7be_uxn_opcodes_h_l1189_c3_f7be_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1193_c11_cac5]
signal BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1193_c7_3e75]
signal t8_MUX_uxn_opcodes_h_l1193_c7_3e75_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1193_c7_3e75]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1193_c7_3e75]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1193_c7_3e75]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1193_c7_3e75]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1193_c7_3e75]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1193_c7_3e75]
signal result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1193_c7_3e75]
signal n8_MUX_uxn_opcodes_h_l1193_c7_3e75_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1196_c11_1c7e]
signal BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1196_c7_dc40]
signal t8_MUX_uxn_opcodes_h_l1196_c7_dc40_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1196_c7_dc40]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1196_c7_dc40]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1196_c7_dc40]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1196_c7_dc40]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1196_c7_dc40]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1196_c7_dc40]
signal result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1196_c7_dc40]
signal n8_MUX_uxn_opcodes_h_l1196_c7_dc40_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1199_c11_24da]
signal BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1199_c7_0ac2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1199_c7_0ac2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1199_c7_0ac2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1199_c7_0ac2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1199_c7_0ac2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1199_c7_0ac2]
signal result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1199_c7_0ac2]
signal n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1202_c30_b18c]
signal sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1205_c21_7e6c]
signal BIN_OP_EQ_uxn_opcodes_h_l1205_c21_7e6c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1205_c21_7e6c_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1205_c21_7e6c_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1205_c21_1654]
signal MUX_uxn_opcodes_h_l1205_c21_1654_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1205_c21_1654_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1205_c21_1654_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1205_c21_1654_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1207_c11_a107]
signal BIN_OP_EQ_uxn_opcodes_h_l1207_c11_a107_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1207_c11_a107_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1207_c11_a107_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1207_c7_d458]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1207_c7_d458]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1207_c7_d458]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8c29( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d
BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_left,
BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_right,
BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_return_output);

-- t8_MUX_uxn_opcodes_h_l1188_c2_5b1f
t8_MUX_uxn_opcodes_h_l1188_c2_5b1f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond,
t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue,
t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse,
t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f
result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f
result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f
result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f
result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output);

-- n8_MUX_uxn_opcodes_h_l1188_c2_5b1f
n8_MUX_uxn_opcodes_h_l1188_c2_5b1f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond,
n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue,
n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse,
n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output);

-- printf_uxn_opcodes_h_l1189_c3_f7be_uxn_opcodes_h_l1189_c3_f7be
printf_uxn_opcodes_h_l1189_c3_f7be_uxn_opcodes_h_l1189_c3_f7be : entity work.printf_uxn_opcodes_h_l1189_c3_f7be_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1189_c3_f7be_uxn_opcodes_h_l1189_c3_f7be_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5
BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_left,
BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_right,
BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_return_output);

-- t8_MUX_uxn_opcodes_h_l1193_c7_3e75
t8_MUX_uxn_opcodes_h_l1193_c7_3e75 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1193_c7_3e75_cond,
t8_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue,
t8_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse,
t8_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75
result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75
result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75
result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75
result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75
result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_cond,
result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output);

-- n8_MUX_uxn_opcodes_h_l1193_c7_3e75
n8_MUX_uxn_opcodes_h_l1193_c7_3e75 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1193_c7_3e75_cond,
n8_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue,
n8_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse,
n8_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e
BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_left,
BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_right,
BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_return_output);

-- t8_MUX_uxn_opcodes_h_l1196_c7_dc40
t8_MUX_uxn_opcodes_h_l1196_c7_dc40 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1196_c7_dc40_cond,
t8_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue,
t8_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse,
t8_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40
result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40
result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40
result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40
result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40
result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_cond,
result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output);

-- n8_MUX_uxn_opcodes_h_l1196_c7_dc40
n8_MUX_uxn_opcodes_h_l1196_c7_dc40 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1196_c7_dc40_cond,
n8_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue,
n8_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse,
n8_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da
BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_left,
BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_right,
BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2
result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2
result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2
result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond,
result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output);

-- n8_MUX_uxn_opcodes_h_l1199_c7_0ac2
n8_MUX_uxn_opcodes_h_l1199_c7_0ac2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond,
n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue,
n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse,
n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c
sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_ins,
sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_x,
sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_y,
sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1205_c21_7e6c
BIN_OP_EQ_uxn_opcodes_h_l1205_c21_7e6c : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1205_c21_7e6c_left,
BIN_OP_EQ_uxn_opcodes_h_l1205_c21_7e6c_right,
BIN_OP_EQ_uxn_opcodes_h_l1205_c21_7e6c_return_output);

-- MUX_uxn_opcodes_h_l1205_c21_1654
MUX_uxn_opcodes_h_l1205_c21_1654 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1205_c21_1654_cond,
MUX_uxn_opcodes_h_l1205_c21_1654_iftrue,
MUX_uxn_opcodes_h_l1205_c21_1654_iffalse,
MUX_uxn_opcodes_h_l1205_c21_1654_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1207_c11_a107
BIN_OP_EQ_uxn_opcodes_h_l1207_c11_a107 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1207_c11_a107_left,
BIN_OP_EQ_uxn_opcodes_h_l1207_c11_a107_right,
BIN_OP_EQ_uxn_opcodes_h_l1207_c11_a107_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458
result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458
result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458
result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_return_output,
 t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output,
 n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_return_output,
 t8_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output,
 n8_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_return_output,
 t8_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output,
 n8_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output,
 n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output,
 sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1205_c21_7e6c_return_output,
 MUX_uxn_opcodes_h_l1205_c21_1654_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1207_c11_a107_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1190_c3_3381 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1189_c3_f7be_uxn_opcodes_h_l1189_c3_f7be_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1193_c7_3e75_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1194_c3_5661 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1193_c7_3e75_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1196_c7_dc40_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1196_c7_dc40_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1204_c3_0c5a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1205_c21_1654_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1205_c21_1654_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1205_c21_1654_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_7e6c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_7e6c_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_7e6c_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1205_c21_1654_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_a107_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_a107_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_a107_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_f168_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_369f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_0f2f_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_aabf_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1199_l1193_l1207_l1196_DUPLICATE_6ce8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1199_l1196_DUPLICATE_cb4e_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l1213_l1184_DUPLICATE_f841_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_right := to_unsigned(3, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1205_c21_1654_iffalse := resize(to_unsigned(1, 1), 8);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_right := to_unsigned(2, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1190_c3_3381 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1190_c3_3381;
     VAR_MUX_uxn_opcodes_h_l1205_c21_1654_iftrue := resize(to_unsigned(0, 1), 8);
     VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1194_c3_5661 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1194_c3_5661;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_a107_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1204_c3_0c5a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1204_c3_0c5a;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_a107_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_7e6c_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_7e6c_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1196_c11_1c7e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_0f2f LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_0f2f_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_aabf LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_aabf_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1199_l1193_l1207_l1196_DUPLICATE_6ce8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1199_l1193_l1207_l1196_DUPLICATE_6ce8_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1193_c11_cac5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_left;
     BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_return_output := BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1199_l1196_DUPLICATE_cb4e LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1199_l1196_DUPLICATE_cb4e_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_f168 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_f168_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1207_c11_a107] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1207_c11_a107_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_a107_left;
     BIN_OP_EQ_uxn_opcodes_h_l1207_c11_a107_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_a107_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_a107_return_output := BIN_OP_EQ_uxn_opcodes_h_l1207_c11_a107_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_369f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_369f_return_output := result.is_stack_write;

     -- sp_relative_shift[uxn_opcodes_h_l1202_c30_b18c] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_ins;
     sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_x;
     sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_return_output := sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1205_c21_7e6c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1205_c21_7e6c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_7e6c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1205_c21_7e6c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_7e6c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_7e6c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1205_c21_7e6c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1199_c11_24da] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_left;
     BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_return_output := BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1188_c6_7c4d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_7c4d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1193_c7_3e75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1193_c7_3e75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_cac5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1196_c7_dc40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1196_c7_dc40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_1c7e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_24da_return_output;
     VAR_MUX_uxn_opcodes_h_l1205_c21_1654_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_7e6c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_a107_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_a107_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_a107_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_0f2f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_0f2f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_0f2f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_0f2f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1199_l1193_l1207_l1196_DUPLICATE_6ce8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1199_l1193_l1207_l1196_DUPLICATE_6ce8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1199_l1193_l1207_l1196_DUPLICATE_6ce8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1199_l1193_l1207_l1196_DUPLICATE_6ce8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_f168_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_f168_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_f168_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_f168_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_369f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_369f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_369f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_369f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1199_l1196_DUPLICATE_cb4e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1199_l1196_DUPLICATE_cb4e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_aabf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_aabf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_aabf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_aabf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_b18c_return_output;
     -- t8_MUX[uxn_opcodes_h_l1196_c7_dc40] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1196_c7_dc40_cond <= VAR_t8_MUX_uxn_opcodes_h_l1196_c7_dc40_cond;
     t8_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue;
     t8_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output := t8_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output;

     -- n8_MUX[uxn_opcodes_h_l1199_c7_0ac2] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond <= VAR_n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond;
     n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue;
     n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output := n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1207_c7_d458] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1188_c1_afa1] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1199_c7_0ac2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output;

     -- MUX[uxn_opcodes_h_l1205_c21_1654] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1205_c21_1654_cond <= VAR_MUX_uxn_opcodes_h_l1205_c21_1654_cond;
     MUX_uxn_opcodes_h_l1205_c21_1654_iftrue <= VAR_MUX_uxn_opcodes_h_l1205_c21_1654_iftrue;
     MUX_uxn_opcodes_h_l1205_c21_1654_iffalse <= VAR_MUX_uxn_opcodes_h_l1205_c21_1654_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1205_c21_1654_return_output := MUX_uxn_opcodes_h_l1205_c21_1654_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1199_c7_0ac2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1207_c7_d458] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1207_c7_d458] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue := VAR_MUX_uxn_opcodes_h_l1205_c21_1654_return_output;
     VAR_printf_uxn_opcodes_h_l1189_c3_f7be_uxn_opcodes_h_l1189_c3_f7be_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_afa1_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_d458_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_d458_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_d458_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output;
     -- printf_uxn_opcodes_h_l1189_c3_f7be[uxn_opcodes_h_l1189_c3_f7be] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1189_c3_f7be_uxn_opcodes_h_l1189_c3_f7be_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1189_c3_f7be_uxn_opcodes_h_l1189_c3_f7be_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_u8_value_MUX[uxn_opcodes_h_l1199_c7_0ac2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output := result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1196_c7_dc40] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1199_c7_0ac2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output;

     -- t8_MUX[uxn_opcodes_h_l1193_c7_3e75] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1193_c7_3e75_cond <= VAR_t8_MUX_uxn_opcodes_h_l1193_c7_3e75_cond;
     t8_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue;
     t8_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output := t8_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1196_c7_dc40] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output;

     -- n8_MUX[uxn_opcodes_h_l1196_c7_dc40] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1196_c7_dc40_cond <= VAR_n8_MUX_uxn_opcodes_h_l1196_c7_dc40_cond;
     n8_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue;
     n8_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output := n8_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1199_c7_0ac2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1199_c7_0ac2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_0ac2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output;
     -- n8_MUX[uxn_opcodes_h_l1193_c7_3e75] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1193_c7_3e75_cond <= VAR_n8_MUX_uxn_opcodes_h_l1193_c7_3e75_cond;
     n8_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue;
     n8_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output := n8_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1193_c7_3e75] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1196_c7_dc40] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output := result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1196_c7_dc40] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1196_c7_dc40] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1193_c7_3e75] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output;

     -- t8_MUX[uxn_opcodes_h_l1188_c2_5b1f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond <= VAR_t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond;
     t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue;
     t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output := t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1196_c7_dc40] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_dc40_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1188_c2_5b1f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1188_c2_5b1f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1193_c7_3e75] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1193_c7_3e75] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1193_c7_3e75] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output := result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output;

     -- n8_MUX[uxn_opcodes_h_l1188_c2_5b1f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond <= VAR_n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond;
     n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue;
     n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output := n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1193_c7_3e75] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_3e75_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1188_c2_5b1f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1188_c2_5b1f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1188_c2_5b1f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1188_c2_5b1f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l1213_l1184_DUPLICATE_f841 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l1213_l1184_DUPLICATE_f841_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8c29(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_5b1f_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l1213_l1184_DUPLICATE_f841_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l1213_l1184_DUPLICATE_f841_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
