-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 47
entity str1_0CLK_faaf4b1a is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end str1_0CLK_faaf4b1a;
architecture arch of str1_0CLK_faaf4b1a is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1604_c6_03cb]
signal BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1604_c1_54c5]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1604_c2_7d96]
signal t8_MUX_uxn_opcodes_h_l1604_c2_7d96_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1604_c2_7d96]
signal n8_MUX_uxn_opcodes_h_l1604_c2_7d96_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1604_c2_7d96]
signal result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1604_c2_7d96]
signal result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1604_c2_7d96]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1604_c2_7d96]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1604_c2_7d96]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1604_c2_7d96]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output : signed(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1604_c2_7d96]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l1605_c3_e571[uxn_opcodes_h_l1605_c3_e571]
signal printf_uxn_opcodes_h_l1605_c3_e571_uxn_opcodes_h_l1605_c3_e571_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1609_c11_4b96]
signal BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1609_c7_2944]
signal t8_MUX_uxn_opcodes_h_l1609_c7_2944_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1609_c7_2944_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1609_c7_2944]
signal n8_MUX_uxn_opcodes_h_l1609_c7_2944_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1609_c7_2944_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1609_c7_2944]
signal result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1609_c7_2944]
signal result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1609_c7_2944]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1609_c7_2944]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1609_c7_2944]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1609_c7_2944]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_return_output : signed(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1609_c7_2944]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1612_c11_bc76]
signal BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1612_c7_d182]
signal t8_MUX_uxn_opcodes_h_l1612_c7_d182_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1612_c7_d182_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1612_c7_d182]
signal n8_MUX_uxn_opcodes_h_l1612_c7_d182_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1612_c7_d182_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1612_c7_d182]
signal result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1612_c7_d182]
signal result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1612_c7_d182]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1612_c7_d182]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1612_c7_d182]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_return_output : signed(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1612_c7_d182]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1615_c11_025b]
signal BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1615_c7_98be]
signal n8_MUX_uxn_opcodes_h_l1615_c7_98be_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1615_c7_98be_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1615_c7_98be]
signal result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1615_c7_98be]
signal result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1615_c7_98be]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1615_c7_98be]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1615_c7_98be]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_return_output : signed(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1615_c7_98be]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1618_c30_8572]
signal sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_return_output : signed(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1620_c22_abf5]
signal BIN_OP_PLUS_uxn_opcodes_h_l1620_c22_abf5_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1620_c22_abf5_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1620_c22_abf5_return_output : signed(17 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1623_c11_a0a3]
signal BIN_OP_EQ_uxn_opcodes_h_l1623_c11_a0a3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1623_c11_a0a3_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1623_c11_a0a3_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1623_c7_960a]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1623_c7_960a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1623_c7_960a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_return_output : unsigned(0 downto 0);

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_c878( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u16_value := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_ram_write := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb
BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_left,
BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_right,
BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_return_output);

-- t8_MUX_uxn_opcodes_h_l1604_c2_7d96
t8_MUX_uxn_opcodes_h_l1604_c2_7d96 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1604_c2_7d96_cond,
t8_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue,
t8_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse,
t8_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output);

-- n8_MUX_uxn_opcodes_h_l1604_c2_7d96
n8_MUX_uxn_opcodes_h_l1604_c2_7d96 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1604_c2_7d96_cond,
n8_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue,
n8_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse,
n8_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96
result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_cond,
result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96
result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_cond,
result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96
result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96
result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96
result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96
result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output);

-- printf_uxn_opcodes_h_l1605_c3_e571_uxn_opcodes_h_l1605_c3_e571
printf_uxn_opcodes_h_l1605_c3_e571_uxn_opcodes_h_l1605_c3_e571 : entity work.printf_uxn_opcodes_h_l1605_c3_e571_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1605_c3_e571_uxn_opcodes_h_l1605_c3_e571_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96
BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_left,
BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_right,
BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_return_output);

-- t8_MUX_uxn_opcodes_h_l1609_c7_2944
t8_MUX_uxn_opcodes_h_l1609_c7_2944 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1609_c7_2944_cond,
t8_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue,
t8_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse,
t8_MUX_uxn_opcodes_h_l1609_c7_2944_return_output);

-- n8_MUX_uxn_opcodes_h_l1609_c7_2944
n8_MUX_uxn_opcodes_h_l1609_c7_2944 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1609_c7_2944_cond,
n8_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue,
n8_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse,
n8_MUX_uxn_opcodes_h_l1609_c7_2944_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944
result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_cond,
result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944
result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_cond,
result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944
result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944
result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944
result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944
result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76
BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_left,
BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_right,
BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_return_output);

-- t8_MUX_uxn_opcodes_h_l1612_c7_d182
t8_MUX_uxn_opcodes_h_l1612_c7_d182 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1612_c7_d182_cond,
t8_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue,
t8_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse,
t8_MUX_uxn_opcodes_h_l1612_c7_d182_return_output);

-- n8_MUX_uxn_opcodes_h_l1612_c7_d182
n8_MUX_uxn_opcodes_h_l1612_c7_d182 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1612_c7_d182_cond,
n8_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue,
n8_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse,
n8_MUX_uxn_opcodes_h_l1612_c7_d182_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182
result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_cond,
result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182
result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_cond,
result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182
result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182
result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182
result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182
result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b
BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_left,
BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_right,
BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_return_output);

-- n8_MUX_uxn_opcodes_h_l1615_c7_98be
n8_MUX_uxn_opcodes_h_l1615_c7_98be : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1615_c7_98be_cond,
n8_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue,
n8_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse,
n8_MUX_uxn_opcodes_h_l1615_c7_98be_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be
result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_cond,
result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be
result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_cond,
result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be
result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be
result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be
result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be
result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1618_c30_8572
sp_relative_shift_uxn_opcodes_h_l1618_c30_8572 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_ins,
sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_x,
sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_y,
sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1620_c22_abf5
BIN_OP_PLUS_uxn_opcodes_h_l1620_c22_abf5 : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1620_c22_abf5_left,
BIN_OP_PLUS_uxn_opcodes_h_l1620_c22_abf5_right,
BIN_OP_PLUS_uxn_opcodes_h_l1620_c22_abf5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1623_c11_a0a3
BIN_OP_EQ_uxn_opcodes_h_l1623_c11_a0a3 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1623_c11_a0a3_left,
BIN_OP_EQ_uxn_opcodes_h_l1623_c11_a0a3_right,
BIN_OP_EQ_uxn_opcodes_h_l1623_c11_a0a3_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a
result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a
result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a
result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_return_output,
 t8_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output,
 n8_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_return_output,
 t8_MUX_uxn_opcodes_h_l1609_c7_2944_return_output,
 n8_MUX_uxn_opcodes_h_l1609_c7_2944_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_return_output,
 t8_MUX_uxn_opcodes_h_l1612_c7_d182_return_output,
 n8_MUX_uxn_opcodes_h_l1612_c7_d182_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_return_output,
 n8_MUX_uxn_opcodes_h_l1615_c7_98be_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_return_output,
 sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1620_c22_abf5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1623_c11_a0a3_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1609_c7_2944_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1604_c2_7d96_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1609_c7_2944_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1604_c2_7d96_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1606_c3_fa18 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1605_c3_e571_uxn_opcodes_h_l1605_c3_e571_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1612_c7_d182_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1609_c7_2944_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1612_c7_d182_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1609_c7_2944_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1610_c3_2e8a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1609_c7_2944_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1612_c7_d182_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1615_c7_98be_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1612_c7_d182_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1615_c7_98be_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l1620_c3_3acb : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1620_c22_abf5_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l1620_c27_048c_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1620_c22_abf5_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1620_c22_abf5_return_output : signed(17 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1623_c11_a0a3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1623_c11_a0a3_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1623_c11_a0a3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1609_l1612_l1604_l1615_DUPLICATE_f741_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1609_l1612_l1604_l1615_DUPLICATE_5d1a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1609_l1623_l1612_l1604_DUPLICATE_e1ac_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1609_l1612_l1604_l1615_DUPLICATE_168b_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1609_l1623_l1612_l1604_DUPLICATE_ea7d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1609_l1623_l1612_l1615_DUPLICATE_af9b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c878_uxn_opcodes_h_l1629_l1600_DUPLICATE_91f9_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_y := resize(to_signed(-2, 3), 4);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1610_c3_2e8a := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1610_c3_2e8a;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1606_c3_fa18 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1606_c3_fa18;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_right := to_unsigned(2, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1623_c11_a0a3_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse := n8;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1620_c22_abf5_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1623_c11_a0a3_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse := t8;
     -- CAST_TO_int8_t[uxn_opcodes_h_l1620_c27_048c] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l1620_c27_048c_return_output := CAST_TO_int8_t_uint8_t(
     t8);

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1609_l1623_l1612_l1615_DUPLICATE_af9b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1609_l1623_l1612_l1615_DUPLICATE_af9b_return_output := result.is_opc_done;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1609_c7_2944] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1609_c7_2944_return_output := result.stack_address_sp_offset;

     -- sp_relative_shift[uxn_opcodes_h_l1618_c30_8572] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_ins;
     sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_x;
     sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_return_output := sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1609_l1623_l1612_l1604_DUPLICATE_ea7d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1609_l1623_l1612_l1604_DUPLICATE_ea7d_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1609_l1612_l1604_l1615_DUPLICATE_5d1a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1609_l1612_l1604_l1615_DUPLICATE_5d1a_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1604_c6_03cb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_left;
     BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_return_output := BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1615_c11_025b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1609_l1612_l1604_l1615_DUPLICATE_168b LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1609_l1612_l1604_l1615_DUPLICATE_168b_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1609_l1612_l1604_l1615_DUPLICATE_f741 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1609_l1612_l1604_l1615_DUPLICATE_f741_return_output := result.u16_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1609_c11_4b96] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_left;
     BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_return_output := BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1612_c11_bc76] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_left;
     BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_return_output := BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1623_c11_a0a3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1623_c11_a0a3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1623_c11_a0a3_left;
     BIN_OP_EQ_uxn_opcodes_h_l1623_c11_a0a3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1623_c11_a0a3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1623_c11_a0a3_return_output := BIN_OP_EQ_uxn_opcodes_h_l1623_c11_a0a3_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1609_l1623_l1612_l1604_DUPLICATE_e1ac LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1609_l1623_l1612_l1604_DUPLICATE_e1ac_return_output := result.is_sp_shift;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1604_c2_7d96_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1604_c2_7d96_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1604_c6_03cb_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1609_c7_2944_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1609_c7_2944_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1609_c11_4b96_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1612_c7_d182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1612_c7_d182_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1612_c11_bc76_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1615_c7_98be_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1615_c11_025b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1623_c11_a0a3_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1623_c11_a0a3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1623_c11_a0a3_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1620_c22_abf5_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l1620_c27_048c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1609_l1612_l1604_l1615_DUPLICATE_168b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1609_l1612_l1604_l1615_DUPLICATE_168b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1609_l1612_l1604_l1615_DUPLICATE_168b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1609_l1612_l1604_l1615_DUPLICATE_168b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1609_l1612_l1604_l1615_DUPLICATE_f741_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1609_l1612_l1604_l1615_DUPLICATE_f741_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1609_l1612_l1604_l1615_DUPLICATE_f741_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1609_l1612_l1604_l1615_DUPLICATE_f741_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1609_l1623_l1612_l1615_DUPLICATE_af9b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1609_l1623_l1612_l1615_DUPLICATE_af9b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1609_l1623_l1612_l1615_DUPLICATE_af9b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1609_l1623_l1612_l1615_DUPLICATE_af9b_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1609_l1623_l1612_l1604_DUPLICATE_ea7d_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1609_l1623_l1612_l1604_DUPLICATE_ea7d_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1609_l1623_l1612_l1604_DUPLICATE_ea7d_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1609_l1623_l1612_l1604_DUPLICATE_ea7d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1609_l1623_l1612_l1604_DUPLICATE_e1ac_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1609_l1623_l1612_l1604_DUPLICATE_e1ac_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1609_l1623_l1612_l1604_DUPLICATE_e1ac_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1609_l1623_l1612_l1604_DUPLICATE_e1ac_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1609_l1612_l1604_l1615_DUPLICATE_5d1a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1609_l1612_l1604_l1615_DUPLICATE_5d1a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1609_l1612_l1604_l1615_DUPLICATE_5d1a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1609_l1612_l1604_l1615_DUPLICATE_5d1a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1609_c7_2944_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1618_c30_8572_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1615_c7_98be] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1604_c1_54c5] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1615_c7_98be] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_return_output := result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1623_c7_960a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1620_c22_abf5] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1620_c22_abf5_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1620_c22_abf5_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1620_c22_abf5_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1620_c22_abf5_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1620_c22_abf5_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1620_c22_abf5_return_output;

     -- n8_MUX[uxn_opcodes_h_l1615_c7_98be] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1615_c7_98be_cond <= VAR_n8_MUX_uxn_opcodes_h_l1615_c7_98be_cond;
     n8_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue;
     n8_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1615_c7_98be_return_output := n8_MUX_uxn_opcodes_h_l1615_c7_98be_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1623_c7_960a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1623_c7_960a] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1609_c7_2944] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_return_output;

     -- t8_MUX[uxn_opcodes_h_l1612_c7_d182] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1612_c7_d182_cond <= VAR_t8_MUX_uxn_opcodes_h_l1612_c7_d182_cond;
     t8_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue;
     t8_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1612_c7_d182_return_output := t8_MUX_uxn_opcodes_h_l1612_c7_d182_return_output;

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l1620_c3_3acb := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1620_c22_abf5_return_output)),16);
     VAR_printf_uxn_opcodes_h_l1605_c3_e571_uxn_opcodes_h_l1605_c3_e571_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1604_c1_54c5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1615_c7_98be_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1623_c7_960a_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1623_c7_960a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1623_c7_960a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1615_c7_98be_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1609_c7_2944_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1615_c7_98be_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1612_c7_d182_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue := VAR_result_u16_value_uxn_opcodes_h_l1620_c3_3acb;
     -- result_u8_value_MUX[uxn_opcodes_h_l1612_c7_d182] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_return_output := result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1604_c2_7d96] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1615_c7_98be] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1615_c7_98be] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_return_output;

     -- t8_MUX[uxn_opcodes_h_l1609_c7_2944] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1609_c7_2944_cond <= VAR_t8_MUX_uxn_opcodes_h_l1609_c7_2944_cond;
     t8_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue;
     t8_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1609_c7_2944_return_output := t8_MUX_uxn_opcodes_h_l1609_c7_2944_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1615_c7_98be] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1615_c7_98be] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_return_output := result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1612_c7_d182] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_return_output;

     -- printf_uxn_opcodes_h_l1605_c3_e571[uxn_opcodes_h_l1605_c3_e571] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1605_c3_e571_uxn_opcodes_h_l1605_c3_e571_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1605_c3_e571_uxn_opcodes_h_l1605_c3_e571_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- n8_MUX[uxn_opcodes_h_l1612_c7_d182] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1612_c7_d182_cond <= VAR_n8_MUX_uxn_opcodes_h_l1612_c7_d182_cond;
     n8_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue;
     n8_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1612_c7_d182_return_output := n8_MUX_uxn_opcodes_h_l1612_c7_d182_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1612_c7_d182_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1615_c7_98be_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1615_c7_98be_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1615_c7_98be_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1612_c7_d182_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1615_c7_98be_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1612_c7_d182_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1609_c7_2944_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1609_c7_2944] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_return_output := result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1612_c7_d182] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_return_output := result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1612_c7_d182] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1609_c7_2944] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_return_output;

     -- n8_MUX[uxn_opcodes_h_l1609_c7_2944] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1609_c7_2944_cond <= VAR_n8_MUX_uxn_opcodes_h_l1609_c7_2944_cond;
     n8_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue;
     n8_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1609_c7_2944_return_output := n8_MUX_uxn_opcodes_h_l1609_c7_2944_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1612_c7_d182] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_return_output;

     -- t8_MUX[uxn_opcodes_h_l1604_c2_7d96] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1604_c2_7d96_cond <= VAR_t8_MUX_uxn_opcodes_h_l1604_c2_7d96_cond;
     t8_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue;
     t8_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output := t8_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1612_c7_d182] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1609_c7_2944_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1612_c7_d182_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1612_c7_d182_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1612_c7_d182_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1609_c7_2944_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1612_c7_d182_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1609_c7_2944_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1609_c7_2944] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_return_output;

     -- n8_MUX[uxn_opcodes_h_l1604_c2_7d96] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1604_c2_7d96_cond <= VAR_n8_MUX_uxn_opcodes_h_l1604_c2_7d96_cond;
     n8_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue;
     n8_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output := n8_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1609_c7_2944] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_return_output := result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1609_c7_2944] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1609_c7_2944] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1604_c2_7d96] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1604_c2_7d96] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output := result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1609_c7_2944_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1609_c7_2944_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1609_c7_2944_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1609_c7_2944_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1604_c2_7d96] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1604_c2_7d96] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1604_c2_7d96] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1604_c2_7d96] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output := result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c878_uxn_opcodes_h_l1629_l1600_DUPLICATE_91f9 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c878_uxn_opcodes_h_l1629_l1600_DUPLICATE_91f9_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c878(
     result,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1604_c2_7d96_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c878_uxn_opcodes_h_l1629_l1600_DUPLICATE_91f9_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c878_uxn_opcodes_h_l1629_l1600_DUPLICATE_91f9_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
