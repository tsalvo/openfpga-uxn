-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity rot_0CLK_b288bfb7 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end rot_0CLK_b288bfb7;
architecture arch of rot_0CLK_b288bfb7 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal l8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_l8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2657_c6_0033]
signal BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2657_c2_03e7]
signal t8_MUX_uxn_opcodes_h_l2657_c2_03e7_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2657_c2_03e7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2657_c2_03e7]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2657_c2_03e7]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2657_c2_03e7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2657_c2_03e7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2657_c2_03e7]
signal result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2657_c2_03e7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2657_c2_03e7]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2657_c2_03e7]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2657_c2_03e7]
signal l8_MUX_uxn_opcodes_h_l2657_c2_03e7_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2657_c2_03e7]
signal n8_MUX_uxn_opcodes_h_l2657_c2_03e7_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2670_c11_de00]
signal BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2670_c7_0ca0]
signal t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2670_c7_0ca0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2670_c7_0ca0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2670_c7_0ca0]
signal result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2670_c7_0ca0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2670_c7_0ca0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output : signed(3 downto 0);

-- l8_MUX[uxn_opcodes_h_l2670_c7_0ca0]
signal l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2670_c7_0ca0]
signal n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2673_c11_36e9]
signal BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2673_c7_b3e0]
signal t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2673_c7_b3e0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2673_c7_b3e0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2673_c7_b3e0]
signal result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2673_c7_b3e0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2673_c7_b3e0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output : signed(3 downto 0);

-- l8_MUX[uxn_opcodes_h_l2673_c7_b3e0]
signal l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2673_c7_b3e0]
signal n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2677_c11_5c8f]
signal BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2677_c7_a66c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2677_c7_a66c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2677_c7_a66c]
signal result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2677_c7_a66c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2677_c7_a66c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output : signed(3 downto 0);

-- l8_MUX[uxn_opcodes_h_l2677_c7_a66c]
signal l8_MUX_uxn_opcodes_h_l2677_c7_a66c_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2677_c7_a66c]
signal n8_MUX_uxn_opcodes_h_l2677_c7_a66c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2679_c30_87f8]
signal sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2684_c11_2be9]
signal BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2684_c7_c384]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2684_c7_c384]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2684_c7_c384]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2684_c7_c384]
signal result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l2684_c7_c384]
signal l8_MUX_uxn_opcodes_h_l2684_c7_c384_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2684_c7_c384_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2690_c11_9c9b]
signal BIN_OP_EQ_uxn_opcodes_h_l2690_c11_9c9b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2690_c11_9c9b_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2690_c11_9c9b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2690_c7_2d3d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2690_c7_2d3d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2690_c7_2d3d]
signal result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c580( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.u8_value := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_stack_index_flipped := ref_toks_8;
      base.is_pc_updated := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033
BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_left,
BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_right,
BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_return_output);

-- t8_MUX_uxn_opcodes_h_l2657_c2_03e7
t8_MUX_uxn_opcodes_h_l2657_c2_03e7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2657_c2_03e7_cond,
t8_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue,
t8_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse,
t8_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7
result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7
result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7
result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7
result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7
result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_cond,
result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7
result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7
result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output);

-- l8_MUX_uxn_opcodes_h_l2657_c2_03e7
l8_MUX_uxn_opcodes_h_l2657_c2_03e7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2657_c2_03e7_cond,
l8_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue,
l8_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse,
l8_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output);

-- n8_MUX_uxn_opcodes_h_l2657_c2_03e7
n8_MUX_uxn_opcodes_h_l2657_c2_03e7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2657_c2_03e7_cond,
n8_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue,
n8_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse,
n8_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00
BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_left,
BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_right,
BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_return_output);

-- t8_MUX_uxn_opcodes_h_l2670_c7_0ca0
t8_MUX_uxn_opcodes_h_l2670_c7_0ca0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond,
t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue,
t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse,
t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0
result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0
result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond,
result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0
result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0
result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output);

-- l8_MUX_uxn_opcodes_h_l2670_c7_0ca0
l8_MUX_uxn_opcodes_h_l2670_c7_0ca0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond,
l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue,
l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse,
l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output);

-- n8_MUX_uxn_opcodes_h_l2670_c7_0ca0
n8_MUX_uxn_opcodes_h_l2670_c7_0ca0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond,
n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue,
n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse,
n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9
BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_left,
BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_right,
BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_return_output);

-- t8_MUX_uxn_opcodes_h_l2673_c7_b3e0
t8_MUX_uxn_opcodes_h_l2673_c7_b3e0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond,
t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue,
t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse,
t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond,
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0
result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0
result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output);

-- l8_MUX_uxn_opcodes_h_l2673_c7_b3e0
l8_MUX_uxn_opcodes_h_l2673_c7_b3e0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond,
l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue,
l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse,
l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output);

-- n8_MUX_uxn_opcodes_h_l2673_c7_b3e0
n8_MUX_uxn_opcodes_h_l2673_c7_b3e0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond,
n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue,
n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse,
n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f
BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_left,
BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_right,
BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c
result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c
result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c
result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output);

-- l8_MUX_uxn_opcodes_h_l2677_c7_a66c
l8_MUX_uxn_opcodes_h_l2677_c7_a66c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2677_c7_a66c_cond,
l8_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue,
l8_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse,
l8_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output);

-- n8_MUX_uxn_opcodes_h_l2677_c7_a66c
n8_MUX_uxn_opcodes_h_l2677_c7_a66c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2677_c7_a66c_cond,
n8_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue,
n8_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse,
n8_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8
sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_ins,
sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_x,
sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_y,
sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9
BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9_left,
BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9_right,
BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384
result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384
result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384
result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_cond,
result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_return_output);

-- l8_MUX_uxn_opcodes_h_l2684_c7_c384
l8_MUX_uxn_opcodes_h_l2684_c7_c384 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2684_c7_c384_cond,
l8_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue,
l8_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse,
l8_MUX_uxn_opcodes_h_l2684_c7_c384_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2690_c11_9c9b
BIN_OP_EQ_uxn_opcodes_h_l2690_c11_9c9b : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2690_c11_9c9b_left,
BIN_OP_EQ_uxn_opcodes_h_l2690_c11_9c9b_right,
BIN_OP_EQ_uxn_opcodes_h_l2690_c11_9c9b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d
result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d
result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_cond,
result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 l8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_return_output,
 t8_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output,
 l8_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output,
 n8_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_return_output,
 t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output,
 l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output,
 n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_return_output,
 t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output,
 l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output,
 n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output,
 l8_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output,
 n8_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output,
 sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_return_output,
 l8_MUX_uxn_opcodes_h_l2684_c7_c384_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2690_c11_9c9b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2657_c2_03e7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2667_c3_b4c1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2662_c3_72cd : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2657_c2_03e7_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2657_c2_03e7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2671_c3_e72f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2674_c3_a5d5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2681_c3_a8ae : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2684_c7_c384_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2677_c7_a66c_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2677_c7_a66c_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2687_c3_1f77 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2686_c3_25fd : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2684_c7_c384_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_9c9b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_9c9b_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_9c9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2691_c3_2376 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2690_c7_2d3d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2673_l2690_l2657_l2670_DUPLICATE_7a8b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2673_l2670_l2690_l2684_l2677_DUPLICATE_4e65_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2673_l2677_l2670_DUPLICATE_5255_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2673_l2670_l2684_DUPLICATE_17b5_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l2696_l2653_DUPLICATE_7e8e_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_l8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_l8 := l8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2662_c3_72cd := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2662_c3_72cd;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2681_c3_a8ae := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2681_c3_a8ae;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_9c9b_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2691_c3_2376 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2691_c3_2376;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2674_c3_a5d5 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2674_c3_a5d5;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2686_c3_25fd := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2686_c3_25fd;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2667_c3_b4c1 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2667_c3_b4c1;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2687_c3_1f77 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2687_c3_1f77;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2671_c3_e72f := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2671_c3_e72f;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_ins := VAR_ins;
     VAR_l8_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse := l8;
     VAR_n8_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_9c9b_left := VAR_phase;
     VAR_l8_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2684_c11_2be9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9_left;
     BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9_return_output := BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2657_c2_03e7] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2657_c2_03e7_return_output := result.is_vram_write;

     -- sp_relative_shift[uxn_opcodes_h_l2679_c30_87f8] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_ins;
     sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_x;
     sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_return_output := sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2657_c6_0033] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_left;
     BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_return_output := BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2673_l2670_l2690_l2684_l2677_DUPLICATE_4e65 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2673_l2670_l2690_l2684_l2677_DUPLICATE_4e65_return_output := result.is_opc_done;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2657_c2_03e7] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2657_c2_03e7_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2670_c11_de00] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_left;
     BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_return_output := BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2673_c11_36e9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_left;
     BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_return_output := BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2657_c2_03e7] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2657_c2_03e7_return_output := result.is_pc_updated;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2673_l2670_l2684_DUPLICATE_17b5 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2673_l2670_l2684_DUPLICATE_17b5_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2677_c11_5c8f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2690_c7_2d3d] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2690_c7_2d3d_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2673_l2677_l2670_DUPLICATE_5255 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2673_l2677_l2670_DUPLICATE_5255_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2690_c11_9c9b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2690_c11_9c9b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_9c9b_left;
     BIN_OP_EQ_uxn_opcodes_h_l2690_c11_9c9b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_9c9b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_9c9b_return_output := BIN_OP_EQ_uxn_opcodes_h_l2690_c11_9c9b_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2657_c2_03e7] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2657_c2_03e7_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2673_l2690_l2657_l2670_DUPLICATE_7a8b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2673_l2690_l2657_l2670_DUPLICATE_7a8b_return_output := result.u8_value;

     -- Submodule level 1
     VAR_l8_MUX_uxn_opcodes_h_l2657_c2_03e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2657_c2_03e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2657_c2_03e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2657_c6_0033_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2670_c11_de00_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_36e9_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2677_c7_a66c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2677_c7_a66c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2677_c11_5c8f_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2684_c7_c384_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2684_c11_2be9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_9c9b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_9c9b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_9c9b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2673_l2670_l2684_DUPLICATE_17b5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2673_l2670_l2684_DUPLICATE_17b5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2673_l2670_l2684_DUPLICATE_17b5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2673_l2670_l2690_l2684_l2677_DUPLICATE_4e65_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2673_l2670_l2690_l2684_l2677_DUPLICATE_4e65_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2673_l2670_l2690_l2684_l2677_DUPLICATE_4e65_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2673_l2670_l2690_l2684_l2677_DUPLICATE_4e65_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2673_l2670_l2690_l2684_l2677_DUPLICATE_4e65_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2673_l2677_l2670_DUPLICATE_5255_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2673_l2677_l2670_DUPLICATE_5255_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2673_l2677_l2670_DUPLICATE_5255_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2673_l2690_l2657_l2670_DUPLICATE_7a8b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2673_l2690_l2657_l2670_DUPLICATE_7a8b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2673_l2690_l2657_l2670_DUPLICATE_7a8b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2673_l2690_l2657_l2670_DUPLICATE_7a8b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2657_c2_03e7_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2657_c2_03e7_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2657_c2_03e7_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2657_c2_03e7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2690_c7_2d3d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2679_c30_87f8_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2690_c7_2d3d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_return_output;

     -- l8_MUX[uxn_opcodes_h_l2684_c7_c384] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2684_c7_c384_cond <= VAR_l8_MUX_uxn_opcodes_h_l2684_c7_c384_cond;
     l8_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue;
     l8_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2684_c7_c384_return_output := l8_MUX_uxn_opcodes_h_l2684_c7_c384_return_output;

     -- n8_MUX[uxn_opcodes_h_l2677_c7_a66c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2677_c7_a66c_cond <= VAR_n8_MUX_uxn_opcodes_h_l2677_c7_a66c_cond;
     n8_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue;
     n8_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output := n8_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2684_c7_c384] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2657_c2_03e7] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2677_c7_a66c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2657_c2_03e7] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2657_c2_03e7] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2690_c7_2d3d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2657_c2_03e7] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output;

     -- t8_MUX[uxn_opcodes_h_l2673_c7_b3e0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond <= VAR_t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond;
     t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue;
     t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output := t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2690_c7_2d3d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_return_output := result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_return_output;

     -- Submodule level 2
     VAR_l8_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2684_c7_c384_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_2d3d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2684_c7_c384_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_2d3d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2690_c7_2d3d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2684_c7_c384] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_return_output := result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_return_output;

     -- t8_MUX[uxn_opcodes_h_l2670_c7_0ca0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond <= VAR_t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond;
     t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue;
     t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output := t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2673_c7_b3e0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output;

     -- l8_MUX[uxn_opcodes_h_l2677_c7_a66c] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2677_c7_a66c_cond <= VAR_l8_MUX_uxn_opcodes_h_l2677_c7_a66c_cond;
     l8_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue;
     l8_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output := l8_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2684_c7_c384] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2684_c7_c384] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2677_c7_a66c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output;

     -- n8_MUX[uxn_opcodes_h_l2673_c7_b3e0] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond <= VAR_n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond;
     n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue;
     n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output := n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output;

     -- Submodule level 3
     VAR_l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2684_c7_c384_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2684_c7_c384_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2684_c7_c384_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2677_c7_a66c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2670_c7_0ca0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2677_c7_a66c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2673_c7_b3e0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output;

     -- l8_MUX[uxn_opcodes_h_l2673_c7_b3e0] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond <= VAR_l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond;
     l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue;
     l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output := l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2677_c7_a66c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output;

     -- n8_MUX[uxn_opcodes_h_l2670_c7_0ca0] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond <= VAR_n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond;
     n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue;
     n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output := n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output;

     -- t8_MUX[uxn_opcodes_h_l2657_c2_03e7] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2657_c2_03e7_cond <= VAR_t8_MUX_uxn_opcodes_h_l2657_c2_03e7_cond;
     t8_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue;
     t8_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output := t8_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output;

     -- Submodule level 4
     VAR_l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2677_c7_a66c_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2673_c7_b3e0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output := result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output;

     -- l8_MUX[uxn_opcodes_h_l2670_c7_0ca0] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond <= VAR_l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond;
     l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue;
     l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output := l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2673_c7_b3e0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2657_c2_03e7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output;

     -- n8_MUX[uxn_opcodes_h_l2657_c2_03e7] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2657_c2_03e7_cond <= VAR_n8_MUX_uxn_opcodes_h_l2657_c2_03e7_cond;
     n8_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue;
     n8_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output := n8_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2670_c7_0ca0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2673_c7_b3e0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output;

     -- Submodule level 5
     VAR_l8_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output;
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_b3e0_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2670_c7_0ca0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2670_c7_0ca0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output := result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2657_c2_03e7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2670_c7_0ca0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output;

     -- l8_MUX[uxn_opcodes_h_l2657_c2_03e7] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2657_c2_03e7_cond <= VAR_l8_MUX_uxn_opcodes_h_l2657_c2_03e7_cond;
     l8_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue;
     l8_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output := l8_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output;

     -- Submodule level 6
     REG_VAR_l8 := VAR_l8_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2670_c7_0ca0_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2657_c2_03e7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2657_c2_03e7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2657_c2_03e7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output := result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l2696_l2653_DUPLICATE_7e8e LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l2696_l2653_DUPLICATE_7e8e_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c580(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2657_c2_03e7_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l2696_l2653_DUPLICATE_7e8e_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l2696_l2653_DUPLICATE_7e8e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_l8 <= REG_VAR_l8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     l8 <= REG_COMB_l8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
