-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 36
entity nip2_0CLK_1a2ef46d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end nip2_0CLK_1a2ef46d;
architecture arch of nip2_0CLK_1a2ef46d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2174_c6_6a19]
signal BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2174_c2_f45f]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2174_c2_f45f]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2174_c2_f45f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2174_c2_f45f]
signal result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2174_c2_f45f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2174_c2_f45f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2174_c2_f45f]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2174_c2_f45f]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2174_c2_f45f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output : unsigned(3 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2174_c2_f45f]
signal t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output : unsigned(7 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2174_c2_f45f]
signal t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2187_c11_9a4d]
signal BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2187_c7_0a4f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2187_c7_0a4f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2187_c7_0a4f]
signal result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2187_c7_0a4f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2187_c7_0a4f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output : unsigned(3 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2187_c7_0a4f]
signal t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output : unsigned(7 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2187_c7_0a4f]
signal t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2190_c11_8f3f]
signal BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2190_c7_9b48]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2190_c7_9b48]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2190_c7_9b48]
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2190_c7_9b48]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2190_c7_9b48]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output : unsigned(3 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2190_c7_9b48]
signal t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output : unsigned(7 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2190_c7_9b48]
signal t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2192_c30_9580]
signal sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2197_c11_7b8a]
signal BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2197_c7_c597]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2197_c7_c597]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2197_c7_c597]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2197_c7_c597]
signal result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_return_output : unsigned(7 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2197_c7_c597]
signal t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_71f0( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_index_flipped := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.stack_address_sp_offset := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19
BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_left,
BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_right,
BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f
result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f
result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f
result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f
result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f
result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f
result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f
t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_cond,
t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue,
t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse,
t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f
t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_cond,
t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue,
t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse,
t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d
BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_left,
BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_right,
BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f
t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond,
t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue,
t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse,
t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f
t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond,
t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue,
t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse,
t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f
BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_left,
BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_right,
BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_cond,
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48
t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_cond,
t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue,
t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse,
t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48
t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_cond,
t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue,
t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse,
t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2192_c30_9580
sp_relative_shift_uxn_opcodes_h_l2192_c30_9580 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_ins,
sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_x,
sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_y,
sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a
BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a_left,
BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a_right,
BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_cond,
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2197_c7_c597
t16_low_MUX_uxn_opcodes_h_l2197_c7_c597 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_cond,
t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue,
t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse,
t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output,
 t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output,
 t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output,
 t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output,
 t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output,
 t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output,
 t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output,
 sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_return_output,
 t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2174_c2_f45f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2174_c2_f45f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2179_c3_7780 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2174_c2_f45f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2174_c2_f45f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2184_c3_2796 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2188_c3_b286 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2194_c3_a54d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2200_c3_22a6 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2197_c7_c597_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2199_c3_adad : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2187_l2174_l2197_DUPLICATE_2ed3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_cc73_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2187_l2197_DUPLICATE_4863_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2187_l2190_l2197_DUPLICATE_eae1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l2205_l2170_DUPLICATE_9ffd_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2199_c3_adad := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2199_c3_adad;
     VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_y := resize(to_signed(-2, 3), 4);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2200_c3_22a6 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2200_c3_22a6;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2188_c3_b286 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2188_c3_b286;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_right := to_unsigned(2, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2179_c3_7780 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2179_c3_7780;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2184_c3_2796 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2184_c3_2796;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2194_c3_a54d := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2194_c3_a54d;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue := VAR_previous_stack_read;
     VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse := t16_high;
     VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse := t16_low;
     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2187_l2197_DUPLICATE_4863 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2187_l2197_DUPLICATE_4863_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2187_c11_9a4d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_left;
     BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_return_output := BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2174_c2_f45f] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2174_c2_f45f_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_cc73 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_cc73_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2187_l2174_l2197_DUPLICATE_2ed3 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2187_l2174_l2197_DUPLICATE_2ed3_return_output := result.u8_value;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2174_c2_f45f] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2174_c2_f45f_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2197_c11_7b8a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2187_l2190_l2197_DUPLICATE_eae1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2187_l2190_l2197_DUPLICATE_eae1_return_output := result.is_opc_done;

     -- sp_relative_shift[uxn_opcodes_h_l2192_c30_9580] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_ins;
     sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_x;
     sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_return_output := sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2197_c7_c597] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2197_c7_c597_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2174_c6_6a19] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_left;
     BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_return_output := BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2174_c2_f45f] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2174_c2_f45f_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l2190_c11_8f3f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2174_c2_f45f] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2174_c2_f45f_return_output := result.is_pc_updated;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_6a19_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_9a4d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_8f3f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_7b8a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2187_l2197_DUPLICATE_4863_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2187_l2197_DUPLICATE_4863_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2187_l2190_l2197_DUPLICATE_eae1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2187_l2190_l2197_DUPLICATE_eae1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2187_l2190_l2197_DUPLICATE_eae1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_cc73_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_cc73_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2187_l2174_l2197_DUPLICATE_2ed3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2187_l2174_l2197_DUPLICATE_2ed3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2187_l2174_l2197_DUPLICATE_2ed3_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2174_c2_f45f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2174_c2_f45f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2174_c2_f45f_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2174_c2_f45f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2197_c7_c597_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_9580_return_output;
     -- t16_low_MUX[uxn_opcodes_h_l2197_c7_c597] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_cond;
     t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_return_output := t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2197_c7_c597] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2174_c2_f45f] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2174_c2_f45f] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2197_c7_c597] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2174_c2_f45f] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2197_c7_c597] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_return_output := result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2190_c7_9b48] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_cond;
     t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output := t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2190_c7_9b48] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2197_c7_c597] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2174_c2_f45f] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_c597_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_c597_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_c597_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_c597_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_c597_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2190_c7_9b48] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output := result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2187_c7_0a4f] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond;
     t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output := t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2187_c7_0a4f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2190_c7_9b48] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2190_c7_9b48] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2190_c7_9b48] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2190_c7_9b48] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_cond;
     t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output := t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_9b48_return_output;
     -- t16_high_MUX[uxn_opcodes_h_l2174_c2_f45f] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_cond;
     t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output := t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2174_c2_f45f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2187_c7_0a4f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2187_c7_0a4f] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond;
     t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output := t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2187_c7_0a4f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2187_c7_0a4f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2187_c7_0a4f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output;
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_0a4f_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2174_c2_f45f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2174_c2_f45f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2174_c2_f45f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2174_c2_f45f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2174_c2_f45f] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_cond;
     t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output := t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output;

     -- Submodule level 5
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l2205_l2170_DUPLICATE_9ffd LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l2205_l2170_DUPLICATE_9ffd_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_71f0(
     result,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f45f_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l2205_l2170_DUPLICATE_9ffd_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l2205_l2170_DUPLICATE_9ffd_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
