-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 46
entity stz_0CLK_ffdfe23b is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end stz_0CLK_ffdfe23b;
architecture arch of stz_0CLK_ffdfe23b is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1449_c6_e0e9]
signal BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1449_c1_d74d]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1449_c2_b2f5]
signal t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1449_c2_b2f5]
signal n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1449_c2_b2f5]
signal result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1449_c2_b2f5]
signal result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1449_c2_b2f5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1449_c2_b2f5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1449_c2_b2f5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1449_c2_b2f5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output : signed(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1449_c2_b2f5]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l1450_c3_f275[uxn_opcodes_h_l1450_c3_f275]
signal printf_uxn_opcodes_h_l1450_c3_f275_uxn_opcodes_h_l1450_c3_f275_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1454_c11_02f1]
signal BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1454_c7_2ae1]
signal t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1454_c7_2ae1]
signal n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1454_c7_2ae1]
signal result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1454_c7_2ae1]
signal result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1454_c7_2ae1]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1454_c7_2ae1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1454_c7_2ae1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1454_c7_2ae1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output : signed(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1454_c7_2ae1]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1457_c11_dbfe]
signal BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1457_c7_6f6b]
signal t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1457_c7_6f6b]
signal n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1457_c7_6f6b]
signal result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1457_c7_6f6b]
signal result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1457_c7_6f6b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1457_c7_6f6b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1457_c7_6f6b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output : signed(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1457_c7_6f6b]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1460_c11_b4aa]
signal BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1460_c7_8731]
signal n8_MUX_uxn_opcodes_h_l1460_c7_8731_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1460_c7_8731_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1460_c7_8731]
signal result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1460_c7_8731]
signal result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1460_c7_8731]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1460_c7_8731]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1460_c7_8731]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_return_output : signed(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1460_c7_8731]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1463_c30_f8b1]
signal sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1468_c11_b336]
signal BIN_OP_EQ_uxn_opcodes_h_l1468_c11_b336_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1468_c11_b336_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1468_c11_b336_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1468_c7_357a]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1468_c7_357a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1468_c7_357a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_return_output : unsigned(0 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_c878( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u16_value := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_ram_write := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9
BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_left,
BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_right,
BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_return_output);

-- t8_MUX_uxn_opcodes_h_l1449_c2_b2f5
t8_MUX_uxn_opcodes_h_l1449_c2_b2f5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond,
t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue,
t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse,
t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output);

-- n8_MUX_uxn_opcodes_h_l1449_c2_b2f5
n8_MUX_uxn_opcodes_h_l1449_c2_b2f5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond,
n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue,
n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse,
n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5
result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond,
result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5
result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond,
result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5
result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5
result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5
result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5
result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output);

-- printf_uxn_opcodes_h_l1450_c3_f275_uxn_opcodes_h_l1450_c3_f275
printf_uxn_opcodes_h_l1450_c3_f275_uxn_opcodes_h_l1450_c3_f275 : entity work.printf_uxn_opcodes_h_l1450_c3_f275_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1450_c3_f275_uxn_opcodes_h_l1450_c3_f275_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1
BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_left,
BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_right,
BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_return_output);

-- t8_MUX_uxn_opcodes_h_l1454_c7_2ae1
t8_MUX_uxn_opcodes_h_l1454_c7_2ae1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond,
t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue,
t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse,
t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output);

-- n8_MUX_uxn_opcodes_h_l1454_c7_2ae1
n8_MUX_uxn_opcodes_h_l1454_c7_2ae1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond,
n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue,
n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse,
n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1
result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond,
result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1
result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond,
result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1
result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1
result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1
result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1
result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe
BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_left,
BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_right,
BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_return_output);

-- t8_MUX_uxn_opcodes_h_l1457_c7_6f6b
t8_MUX_uxn_opcodes_h_l1457_c7_6f6b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond,
t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue,
t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse,
t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output);

-- n8_MUX_uxn_opcodes_h_l1457_c7_6f6b
n8_MUX_uxn_opcodes_h_l1457_c7_6f6b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond,
n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue,
n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse,
n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b
result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond,
result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b
result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b
result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b
result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b
result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa
BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_left,
BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_right,
BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_return_output);

-- n8_MUX_uxn_opcodes_h_l1460_c7_8731
n8_MUX_uxn_opcodes_h_l1460_c7_8731 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1460_c7_8731_cond,
n8_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue,
n8_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse,
n8_MUX_uxn_opcodes_h_l1460_c7_8731_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731
result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_cond,
result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731
result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_cond,
result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731
result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731
result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731
result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731
result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1
sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_ins,
sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_x,
sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_y,
sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1468_c11_b336
BIN_OP_EQ_uxn_opcodes_h_l1468_c11_b336 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1468_c11_b336_left,
BIN_OP_EQ_uxn_opcodes_h_l1468_c11_b336_right,
BIN_OP_EQ_uxn_opcodes_h_l1468_c11_b336_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a
result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a
result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a
result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_return_output,
 t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output,
 n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_return_output,
 t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output,
 n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_return_output,
 t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output,
 n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_return_output,
 n8_MUX_uxn_opcodes_h_l1460_c7_8731_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_return_output,
 sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1468_c11_b336_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1451_c3_ad8f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1450_c3_f275_uxn_opcodes_h_l1450_c3_f275_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1455_c3_a8d2 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1454_c7_2ae1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1460_c7_8731_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1460_c7_8731_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1465_c22_5883_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1468_c11_b336_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1468_c11_b336_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1468_c11_b336_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1449_l1460_l1454_l1457_DUPLICATE_4276_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1449_l1460_l1454_l1457_DUPLICATE_4366_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1449_l1454_l1468_l1457_DUPLICATE_06de_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1449_l1460_l1454_l1457_DUPLICATE_ddfe_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1449_l1454_l1468_l1457_DUPLICATE_1246_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1460_l1454_l1468_l1457_DUPLICATE_12b3_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c878_uxn_opcodes_h_l1474_l1445_DUPLICATE_95f2_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_right := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1451_c3_ad8f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1451_c3_ad8f;
     VAR_sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_y := resize(to_signed(-2, 3), 4);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1455_c3_a8d2 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1455_c3_a8d2;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1468_c11_b336_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_right := to_unsigned(3, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1468_c11_b336_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse := t8;
     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1449_l1460_l1454_l1457_DUPLICATE_ddfe LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1449_l1460_l1454_l1457_DUPLICATE_ddfe_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1449_c6_e0e9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_left;
     BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_return_output := BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1463_c30_f8b1] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_ins;
     sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_x;
     sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_return_output := sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1454_c11_02f1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_left;
     BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_return_output := BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1449_l1454_l1468_l1457_DUPLICATE_06de LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1449_l1454_l1468_l1457_DUPLICATE_06de_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1460_l1454_l1468_l1457_DUPLICATE_12b3 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1460_l1454_l1468_l1457_DUPLICATE_12b3_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1449_l1460_l1454_l1457_DUPLICATE_4366 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1449_l1460_l1454_l1457_DUPLICATE_4366_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1449_l1454_l1468_l1457_DUPLICATE_1246 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1449_l1454_l1468_l1457_DUPLICATE_1246_return_output := result.is_ram_write;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1454_c7_2ae1] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1454_c7_2ae1_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1457_c11_dbfe] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_left;
     BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_return_output := BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_return_output;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1465_c22_5883] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1465_c22_5883_return_output := CAST_TO_uint16_t_uint8_t(
     t8);

     -- BIN_OP_EQ[uxn_opcodes_h_l1460_c11_b4aa] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_left;
     BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_return_output := BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1468_c11_b336] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1468_c11_b336_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1468_c11_b336_left;
     BIN_OP_EQ_uxn_opcodes_h_l1468_c11_b336_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1468_c11_b336_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1468_c11_b336_return_output := BIN_OP_EQ_uxn_opcodes_h_l1468_c11_b336_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1449_l1460_l1454_l1457_DUPLICATE_4276 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1449_l1460_l1454_l1457_DUPLICATE_4276_return_output := result.u16_value;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1449_c6_e0e9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c11_02f1_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1457_c11_dbfe_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1460_c7_8731_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1460_c11_b4aa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1468_c11_b336_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1468_c11_b336_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1468_c11_b336_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1465_c22_5883_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1449_l1460_l1454_l1457_DUPLICATE_ddfe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1449_l1460_l1454_l1457_DUPLICATE_ddfe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1449_l1460_l1454_l1457_DUPLICATE_ddfe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1449_l1460_l1454_l1457_DUPLICATE_ddfe_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1449_l1460_l1454_l1457_DUPLICATE_4276_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1449_l1460_l1454_l1457_DUPLICATE_4276_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1449_l1460_l1454_l1457_DUPLICATE_4276_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1449_l1460_l1454_l1457_DUPLICATE_4276_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1460_l1454_l1468_l1457_DUPLICATE_12b3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1460_l1454_l1468_l1457_DUPLICATE_12b3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1460_l1454_l1468_l1457_DUPLICATE_12b3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1460_l1454_l1468_l1457_DUPLICATE_12b3_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1449_l1454_l1468_l1457_DUPLICATE_1246_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1449_l1454_l1468_l1457_DUPLICATE_1246_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1449_l1454_l1468_l1457_DUPLICATE_1246_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1449_l1454_l1468_l1457_DUPLICATE_1246_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1449_l1454_l1468_l1457_DUPLICATE_06de_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1449_l1454_l1468_l1457_DUPLICATE_06de_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1449_l1454_l1468_l1457_DUPLICATE_06de_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1449_l1454_l1468_l1457_DUPLICATE_06de_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1449_l1460_l1454_l1457_DUPLICATE_4366_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1449_l1460_l1454_l1457_DUPLICATE_4366_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1449_l1460_l1454_l1457_DUPLICATE_4366_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1449_l1460_l1454_l1457_DUPLICATE_4366_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1454_c7_2ae1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1463_c30_f8b1_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1468_c7_357a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_return_output;

     -- t8_MUX[uxn_opcodes_h_l1457_c7_6f6b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond <= VAR_t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond;
     t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue;
     t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output := t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1449_c1_d74d] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1468_c7_357a] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1460_c7_8731] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_return_output := result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_return_output;

     -- n8_MUX[uxn_opcodes_h_l1460_c7_8731] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1460_c7_8731_cond <= VAR_n8_MUX_uxn_opcodes_h_l1460_c7_8731_cond;
     n8_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue;
     n8_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1460_c7_8731_return_output := n8_MUX_uxn_opcodes_h_l1460_c7_8731_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1454_c7_2ae1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1460_c7_8731] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1460_c7_8731] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_return_output := result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1468_c7_357a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l1450_c3_f275_uxn_opcodes_h_l1450_c3_f275_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1449_c1_d74d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1460_c7_8731_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1468_c7_357a_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1468_c7_357a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1468_c7_357a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1460_c7_8731_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1460_c7_8731_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1460_c7_8731_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l1457_c7_6f6b] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output := result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1460_c7_8731] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1460_c7_8731] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_return_output;

     -- printf_uxn_opcodes_h_l1450_c3_f275[uxn_opcodes_h_l1450_c3_f275] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1450_c3_f275_uxn_opcodes_h_l1450_c3_f275_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1450_c3_f275_uxn_opcodes_h_l1450_c3_f275_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- n8_MUX[uxn_opcodes_h_l1457_c7_6f6b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond <= VAR_n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond;
     n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue;
     n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output := n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output;

     -- t8_MUX[uxn_opcodes_h_l1454_c7_2ae1] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond <= VAR_t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond;
     t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue;
     t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output := t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1449_c2_b2f5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1460_c7_8731] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1457_c7_6f6b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1457_c7_6f6b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1460_c7_8731_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1460_c7_8731_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1460_c7_8731_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output;
     -- result_is_ram_write_MUX[uxn_opcodes_h_l1457_c7_6f6b] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1454_c7_2ae1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1454_c7_2ae1] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output := result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output;

     -- n8_MUX[uxn_opcodes_h_l1454_c7_2ae1] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond <= VAR_n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond;
     n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue;
     n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output := n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1457_c7_6f6b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1457_c7_6f6b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output;

     -- t8_MUX[uxn_opcodes_h_l1449_c2_b2f5] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond <= VAR_t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond;
     t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue;
     t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output := t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1454_c7_2ae1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output := result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1457_c7_6f6b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output;
     -- n8_MUX[uxn_opcodes_h_l1449_c2_b2f5] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond <= VAR_n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond;
     n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue;
     n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output := n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1449_c2_b2f5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1449_c2_b2f5] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output := result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1454_c7_2ae1] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1454_c7_2ae1] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1449_c2_b2f5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output := result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1454_c7_2ae1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1454_c7_2ae1_return_output;
     -- result_is_ram_write_MUX[uxn_opcodes_h_l1449_c2_b2f5] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1449_c2_b2f5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1449_c2_b2f5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c878_uxn_opcodes_h_l1474_l1445_DUPLICATE_95f2 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c878_uxn_opcodes_h_l1474_l1445_DUPLICATE_95f2_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c878(
     result,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1449_c2_b2f5_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c878_uxn_opcodes_h_l1474_l1445_DUPLICATE_95f2_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c878_uxn_opcodes_h_l1474_l1445_DUPLICATE_95f2_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
