-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity swp2_0CLK_85d5529e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(15 downto 0);
 return_output : out opcode_result_t);
end swp2_0CLK_85d5529e;
architecture arch of swp2_0CLK_85d5529e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2322_c6_07ca]
signal BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2322_c2_186a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2322_c2_186a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2322_c2_186a]
signal result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2322_c2_186a]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2322_c2_186a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2322_c2_186a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2322_c2_186a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l2322_c2_186a]
signal n16_MUX_uxn_opcodes_h_l2322_c2_186a_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2322_c2_186a_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l2322_c2_186a]
signal t16_MUX_uxn_opcodes_h_l2322_c2_186a_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2322_c2_186a_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2330_c11_b9ed]
signal BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2330_c7_bbd0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2330_c7_bbd0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2330_c7_bbd0]
signal result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2330_c7_bbd0]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2330_c7_bbd0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2330_c7_bbd0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2330_c7_bbd0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l2330_c7_bbd0]
signal n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l2330_c7_bbd0]
signal t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2333_c11_ecfd]
signal BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2333_c7_bdbd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2333_c7_bdbd]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2333_c7_bdbd]
signal result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2333_c7_bdbd]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2333_c7_bdbd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2333_c7_bdbd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2333_c7_bdbd]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l2333_c7_bdbd]
signal n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l2333_c7_bdbd]
signal t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2336_c30_b399]
signal sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2341_c11_4f33]
signal BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2341_c7_4520]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2341_c7_4520]
signal result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2341_c7_4520]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2341_c7_4520]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2341_c7_4520]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2341_c7_4520]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_return_output : unsigned(3 downto 0);

-- n16_MUX[uxn_opcodes_h_l2341_c7_4520]
signal n16_MUX_uxn_opcodes_h_l2341_c7_4520_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l2341_c7_4520_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2347_c11_0c7d]
signal BIN_OP_EQ_uxn_opcodes_h_l2347_c11_0c7d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2347_c11_0c7d_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2347_c11_0c7d_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2347_c7_567c]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2347_c7_567c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2347_c7_567c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8152( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_stack_operation_16bit := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_stack_write := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca
BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_left,
BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_right,
BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a
result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a
result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_cond,
result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a
result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a
result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a
result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_return_output);

-- n16_MUX_uxn_opcodes_h_l2322_c2_186a
n16_MUX_uxn_opcodes_h_l2322_c2_186a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l2322_c2_186a_cond,
n16_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue,
n16_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse,
n16_MUX_uxn_opcodes_h_l2322_c2_186a_return_output);

-- t16_MUX_uxn_opcodes_h_l2322_c2_186a
t16_MUX_uxn_opcodes_h_l2322_c2_186a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2322_c2_186a_cond,
t16_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue,
t16_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse,
t16_MUX_uxn_opcodes_h_l2322_c2_186a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed
BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_left,
BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_right,
BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0
result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0
result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond,
result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0
result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0
result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0
result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output);

-- n16_MUX_uxn_opcodes_h_l2330_c7_bbd0
n16_MUX_uxn_opcodes_h_l2330_c7_bbd0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond,
n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue,
n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse,
n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output);

-- t16_MUX_uxn_opcodes_h_l2330_c7_bbd0
t16_MUX_uxn_opcodes_h_l2330_c7_bbd0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond,
t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue,
t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse,
t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd
BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_left,
BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_right,
BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd
result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd
result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond,
result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd
result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd
result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd
result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output);

-- n16_MUX_uxn_opcodes_h_l2333_c7_bdbd
n16_MUX_uxn_opcodes_h_l2333_c7_bdbd : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond,
n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue,
n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse,
n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output);

-- t16_MUX_uxn_opcodes_h_l2333_c7_bdbd
t16_MUX_uxn_opcodes_h_l2333_c7_bdbd : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond,
t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue,
t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse,
t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2336_c30_b399
sp_relative_shift_uxn_opcodes_h_l2336_c30_b399 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_ins,
sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_x,
sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_y,
sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33
BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_left,
BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_right,
BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520
result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520
result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_cond,
result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520
result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520
result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_return_output);

-- n16_MUX_uxn_opcodes_h_l2341_c7_4520
n16_MUX_uxn_opcodes_h_l2341_c7_4520 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l2341_c7_4520_cond,
n16_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue,
n16_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse,
n16_MUX_uxn_opcodes_h_l2341_c7_4520_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2347_c11_0c7d
BIN_OP_EQ_uxn_opcodes_h_l2347_c11_0c7d : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2347_c11_0c7d_left,
BIN_OP_EQ_uxn_opcodes_h_l2347_c11_0c7d_right,
BIN_OP_EQ_uxn_opcodes_h_l2347_c11_0c7d_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c
result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c
result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_return_output,
 n16_MUX_uxn_opcodes_h_l2322_c2_186a_return_output,
 t16_MUX_uxn_opcodes_h_l2322_c2_186a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output,
 n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output,
 t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output,
 n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output,
 t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output,
 sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_return_output,
 n16_MUX_uxn_opcodes_h_l2341_c7_4520_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2347_c11_0c7d_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2327_c3_07b7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2322_c2_186a_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2322_c2_186a_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2322_c2_186a_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2322_c2_186a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2331_c3_c532 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2338_c3_8b20 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2341_c7_4520_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2344_c3_4b0c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2341_c7_4520_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l2341_c7_4520_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_0c7d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_0c7d_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_0c7d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2341_l2330_l2322_DUPLICATE_811c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2341_l2330_l2322_DUPLICATE_4200_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2330_l2333_l2322_DUPLICATE_d491_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2341_l2330_l2347_l2322_DUPLICATE_034c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2341_l2330_l2347_l2333_DUPLICATE_80ba_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2341_l2330_l2347_l2333_DUPLICATE_4cd0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2353_l2318_DUPLICATE_7c1f_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n16 := n16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2331_c3_c532 := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2331_c3_c532;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2338_c3_8b20 := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2338_c3_8b20;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_0c7d_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2327_c3_07b7 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2327_c3_07b7;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2344_c3_4b0c := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2344_c3_4b0c;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_ins := VAR_ins;
     VAR_n16_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse := n16;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_0c7d_left := VAR_phase;
     VAR_n16_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue := VAR_previous_stack_read;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue := VAR_previous_stack_read;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue := VAR_previous_stack_read;
     VAR_t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue := VAR_previous_stack_read;
     VAR_t16_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse := t16;
     -- BIN_OP_EQ[uxn_opcodes_h_l2347_c11_0c7d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2347_c11_0c7d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_0c7d_left;
     BIN_OP_EQ_uxn_opcodes_h_l2347_c11_0c7d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_0c7d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_0c7d_return_output := BIN_OP_EQ_uxn_opcodes_h_l2347_c11_0c7d_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2330_l2333_l2322_DUPLICATE_d491 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2330_l2333_l2322_DUPLICATE_d491_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2341_l2330_l2347_l2333_DUPLICATE_80ba LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2341_l2330_l2347_l2333_DUPLICATE_80ba_return_output := result.is_stack_operation_16bit;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2341_l2330_l2322_DUPLICATE_4200 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2341_l2330_l2322_DUPLICATE_4200_return_output := result.u16_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2341_c11_4f33] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_left;
     BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_return_output := BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2330_c11_b9ed] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_left;
     BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_return_output := BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2341_l2330_l2347_l2322_DUPLICATE_034c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2341_l2330_l2347_l2322_DUPLICATE_034c_return_output := result.is_stack_write;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2341_c7_4520] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2341_c7_4520_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2341_l2330_l2322_DUPLICATE_811c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2341_l2330_l2322_DUPLICATE_811c_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2341_l2330_l2347_l2333_DUPLICATE_4cd0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2341_l2330_l2347_l2333_DUPLICATE_4cd0_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2322_c6_07ca] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_left;
     BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_return_output := BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2336_c30_b399] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_ins;
     sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_x;
     sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_return_output := sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2333_c11_ecfd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_left;
     BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_return_output := BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_return_output;

     -- Submodule level 1
     VAR_n16_MUX_uxn_opcodes_h_l2322_c2_186a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2322_c2_186a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c6_07ca_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2330_c11_b9ed_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c11_ecfd_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l2341_c7_4520_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_4f33_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_0c7d_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_0c7d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2347_c11_0c7d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2330_l2333_l2322_DUPLICATE_d491_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2330_l2333_l2322_DUPLICATE_d491_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2330_l2333_l2322_DUPLICATE_d491_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2341_l2330_l2322_DUPLICATE_4200_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2341_l2330_l2322_DUPLICATE_4200_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2341_l2330_l2322_DUPLICATE_4200_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2341_l2330_l2347_l2333_DUPLICATE_4cd0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2341_l2330_l2347_l2333_DUPLICATE_4cd0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2341_l2330_l2347_l2333_DUPLICATE_4cd0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2341_l2330_l2347_l2333_DUPLICATE_4cd0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2341_l2330_l2322_DUPLICATE_811c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2341_l2330_l2322_DUPLICATE_811c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2341_l2330_l2322_DUPLICATE_811c_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2341_l2330_l2347_l2333_DUPLICATE_80ba_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2341_l2330_l2347_l2333_DUPLICATE_80ba_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2341_l2330_l2347_l2333_DUPLICATE_80ba_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2341_l2330_l2347_l2333_DUPLICATE_80ba_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2341_l2330_l2347_l2322_DUPLICATE_034c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2341_l2330_l2347_l2322_DUPLICATE_034c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2341_l2330_l2347_l2322_DUPLICATE_034c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2341_l2330_l2347_l2322_DUPLICATE_034c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2341_c7_4520_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2336_c30_b399_return_output;
     -- n16_MUX[uxn_opcodes_h_l2341_c7_4520] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l2341_c7_4520_cond <= VAR_n16_MUX_uxn_opcodes_h_l2341_c7_4520_cond;
     n16_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue;
     n16_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l2341_c7_4520_return_output := n16_MUX_uxn_opcodes_h_l2341_c7_4520_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2341_c7_4520] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2341_c7_4520] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_return_output := result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2347_c7_567c] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2347_c7_567c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2341_c7_4520] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2347_c7_567c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2333_c7_bdbd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output;

     -- t16_MUX[uxn_opcodes_h_l2333_c7_bdbd] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond <= VAR_t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond;
     t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue;
     t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output := t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output;

     -- Submodule level 2
     VAR_n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse := VAR_n16_MUX_uxn_opcodes_h_l2341_c7_4520_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2347_c7_567c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_4520_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2347_c7_567c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2347_c7_567c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_4520_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2341_c7_4520_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2333_c7_bdbd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output;

     -- n16_MUX[uxn_opcodes_h_l2333_c7_bdbd] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond <= VAR_n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond;
     n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue;
     n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output := n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2341_c7_4520] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2333_c7_bdbd] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output := result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2341_c7_4520] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2330_c7_bbd0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output;

     -- t16_MUX[uxn_opcodes_h_l2330_c7_bbd0] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond <= VAR_t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond;
     t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue;
     t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output := t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2341_c7_4520] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2333_c7_bdbd] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output;

     -- Submodule level 3
     VAR_n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse := VAR_n16_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_4520_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2341_c7_4520_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_4520_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2333_c7_bdbd] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2322_c2_186a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_return_output;

     -- n16_MUX[uxn_opcodes_h_l2330_c7_bbd0] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond <= VAR_n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond;
     n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue;
     n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output := n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2330_c7_bbd0] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output := result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2330_c7_bbd0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2333_c7_bdbd] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2333_c7_bdbd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2330_c7_bbd0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output;

     -- t16_MUX[uxn_opcodes_h_l2322_c2_186a] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2322_c2_186a_cond <= VAR_t16_MUX_uxn_opcodes_h_l2322_c2_186a_cond;
     t16_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue;
     t16_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2322_c2_186a_return_output := t16_MUX_uxn_opcodes_h_l2322_c2_186a_return_output;

     -- Submodule level 4
     VAR_n16_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse := VAR_n16_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2333_c7_bdbd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l2322_c2_186a_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2322_c2_186a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2322_c2_186a] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_return_output := result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_return_output;

     -- n16_MUX[uxn_opcodes_h_l2322_c2_186a] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l2322_c2_186a_cond <= VAR_n16_MUX_uxn_opcodes_h_l2322_c2_186a_cond;
     n16_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue;
     n16_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l2322_c2_186a_return_output := n16_MUX_uxn_opcodes_h_l2322_c2_186a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2330_c7_bbd0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2330_c7_bbd0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2330_c7_bbd0] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2322_c2_186a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_return_output;

     -- Submodule level 5
     REG_VAR_n16 := VAR_n16_MUX_uxn_opcodes_h_l2322_c2_186a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2330_c7_bbd0_return_output;
     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2322_c2_186a] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2322_c2_186a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2322_c2_186a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2353_l2318_DUPLICATE_7c1f LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2353_l2318_DUPLICATE_7c1f_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8152(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2322_c2_186a_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2322_c2_186a_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2322_c2_186a_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2322_c2_186a_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2322_c2_186a_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c2_186a_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2322_c2_186a_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2353_l2318_DUPLICATE_7c1f_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l2353_l2318_DUPLICATE_7c1f_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n16 <= REG_VAR_n16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n16 <= REG_COMB_n16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
