-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 49
entity dei_0CLK_9bcaee2f is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_device_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dei_0CLK_9bcaee2f;
architecture arch of dei_0CLK_9bcaee2f is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal has_written_to_t : unsigned(0 downto 0) := to_unsigned(0, 1);
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal device_in_result : device_in_result_t := device_in_result_t_NULL;
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_has_written_to_t : unsigned(0 downto 0);
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_device_in_result : device_in_result_t;
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l403_c6_2848]
signal BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l419_c7_e8d9]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output : unsigned(0 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l403_c2_b756]
signal has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(0 downto 0);

-- device_in_result_MUX[uxn_opcodes_h_l403_c2_b756]
signal device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
signal device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_return_output : device_in_result_t;

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l403_c2_b756]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l403_c2_b756]
signal result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(7 downto 0);

-- result_is_device_ram_write_MUX[uxn_opcodes_h_l403_c2_b756]
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l403_c2_b756]
signal result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l403_c2_b756]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l403_c2_b756]
signal result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l403_c2_b756]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_return_output : signed(3 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l403_c2_b756]
signal result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(7 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l403_c2_b756]
signal result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l403_c2_b756]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l403_c2_b756]
signal result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l403_c2_b756]
signal t8_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l419_c11_29ea]
signal BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l422_c1_340c]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_return_output : unsigned(0 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l419_c7_e8d9]
signal has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output : unsigned(0 downto 0);

-- device_in_result_MUX[uxn_opcodes_h_l419_c7_e8d9]
signal device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_cond : unsigned(0 downto 0);
signal device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output : device_in_result_t;

-- result_device_ram_address_MUX[uxn_opcodes_h_l419_c7_e8d9]
signal result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l419_c7_e8d9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l419_c7_e8d9]
signal result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l419_c7_e8d9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l419_c7_e8d9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l419_c7_e8d9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l419_c7_e8d9]
signal t8_MUX_uxn_opcodes_h_l419_c7_e8d9_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l420_c30_0a72]
signal sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l424_c9_dde0]
signal BIN_OP_EQ_uxn_opcodes_h_l424_c9_dde0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l424_c9_dde0_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l424_c9_dde0_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l424_c9_6298]
signal MUX_uxn_opcodes_h_l424_c9_6298_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l424_c9_6298_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l424_c9_6298_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l424_c9_6298_return_output : unsigned(7 downto 0);

-- UNARY_OP_NOT[uxn_opcodes_h_l425_c8_8f5f]
signal UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8f5f_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8f5f_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l425_c1_46c8]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_return_output : unsigned(0 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l425_c3_8930]
signal has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_return_output : unsigned(0 downto 0);

-- device_in_result_MUX[uxn_opcodes_h_l425_c3_8930]
signal device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_cond : unsigned(0 downto 0);
signal device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_iftrue : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_iffalse : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_return_output : device_in_result_t;

-- result_device_ram_address_MUX[uxn_opcodes_h_l425_c3_8930]
signal result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l425_c3_8930]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l425_c3_8930]
signal result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l425_c3_8930]
signal result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l425_c3_8930]
signal result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_return_output : unsigned(0 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_h_l426_c37_889a]
signal BIN_OP_MINUS_uxn_opcodes_h_l426_c37_889a_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l426_c37_889a_right : unsigned(1 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l426_c37_889a_return_output : unsigned(7 downto 0);

-- device_in[uxn_opcodes_h_l426_c23_b350]
signal device_in_uxn_opcodes_h_l426_c23_b350_CLOCK_ENABLE : unsigned(0 downto 0);
signal device_in_uxn_opcodes_h_l426_c23_b350_device_address : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l426_c23_b350_phase : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l426_c23_b350_previous_device_ram_read : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l426_c23_b350_return_output : device_in_result_t;

-- UNARY_OP_NOT[uxn_opcodes_h_l429_c9_2186]
signal UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2186_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2186_return_output : unsigned(0 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l429_c4_e1db]
signal has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l429_c4_e1db]
signal result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l429_c4_e1db]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l429_c4_e1db]
signal result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l429_c4_e1db]
signal result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_return_output : unsigned(0 downto 0);

function CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6( ref_toks_0 : device_in_result_t;
 ref_toks_1 : unsigned) return device_in_result_t is
 
  variable base : device_in_result_t; 
  variable return_output : device_in_result_t;
begin
      base := ref_toks_0;
      base.is_dei_done := ref_toks_1;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_8fbf( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_device_ram_write := ref_toks_3;
      base.is_ram_write := ref_toks_4;
      base.is_stack_index_flipped := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.device_ram_address := ref_toks_8;
      base.is_vram_write := ref_toks_9;
      base.is_pc_updated := ref_toks_10;
      base.is_opc_done := ref_toks_11;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848
BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_left,
BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_right,
BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_cond,
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_return_output);

-- device_in_result_MUX_uxn_opcodes_h_l403_c2_b756
device_in_result_MUX_uxn_opcodes_h_l403_c2_b756 : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_cond,
device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_iftrue,
device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_iffalse,
device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756
result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_cond,
result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_return_output);

-- result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_cond,
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_iftrue,
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_iffalse,
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_return_output);

-- t8_MUX_uxn_opcodes_h_l403_c2_b756
t8_MUX_uxn_opcodes_h_l403_c2_b756 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l403_c2_b756_cond,
t8_MUX_uxn_opcodes_h_l403_c2_b756_iftrue,
t8_MUX_uxn_opcodes_h_l403_c2_b756_iffalse,
t8_MUX_uxn_opcodes_h_l403_c2_b756_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea
BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_left,
BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_right,
BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_cond,
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output);

-- device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9
device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9 : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_cond,
device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue,
device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse,
device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9
result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_cond,
result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output);

-- t8_MUX_uxn_opcodes_h_l419_c7_e8d9
t8_MUX_uxn_opcodes_h_l419_c7_e8d9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l419_c7_e8d9_cond,
t8_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue,
t8_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse,
t8_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output);

-- sp_relative_shift_uxn_opcodes_h_l420_c30_0a72
sp_relative_shift_uxn_opcodes_h_l420_c30_0a72 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_ins,
sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_x,
sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_y,
sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l424_c9_dde0
BIN_OP_EQ_uxn_opcodes_h_l424_c9_dde0 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l424_c9_dde0_left,
BIN_OP_EQ_uxn_opcodes_h_l424_c9_dde0_right,
BIN_OP_EQ_uxn_opcodes_h_l424_c9_dde0_return_output);

-- MUX_uxn_opcodes_h_l424_c9_6298
MUX_uxn_opcodes_h_l424_c9_6298 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l424_c9_6298_cond,
MUX_uxn_opcodes_h_l424_c9_6298_iftrue,
MUX_uxn_opcodes_h_l424_c9_6298_iffalse,
MUX_uxn_opcodes_h_l424_c9_6298_return_output);

-- UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8f5f
UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8f5f : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8f5f_expr,
UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8f5f_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_cond,
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_return_output);

-- device_in_result_MUX_uxn_opcodes_h_l425_c3_8930
device_in_result_MUX_uxn_opcodes_h_l425_c3_8930 : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_cond,
device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_iftrue,
device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_iffalse,
device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930
result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_cond,
result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l426_c37_889a
BIN_OP_MINUS_uxn_opcodes_h_l426_c37_889a : entity work.BIN_OP_MINUS_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l426_c37_889a_left,
BIN_OP_MINUS_uxn_opcodes_h_l426_c37_889a_right,
BIN_OP_MINUS_uxn_opcodes_h_l426_c37_889a_return_output);

-- device_in_uxn_opcodes_h_l426_c23_b350
device_in_uxn_opcodes_h_l426_c23_b350 : entity work.device_in_0CLK_c6b159da port map (
clk,
device_in_uxn_opcodes_h_l426_c23_b350_CLOCK_ENABLE,
device_in_uxn_opcodes_h_l426_c23_b350_device_address,
device_in_uxn_opcodes_h_l426_c23_b350_phase,
device_in_uxn_opcodes_h_l426_c23_b350_previous_device_ram_read,
device_in_uxn_opcodes_h_l426_c23_b350_return_output);

-- UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2186
UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2186 : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2186_expr,
UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2186_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_cond,
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db
result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_cond,
result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_device_ram_read,
 -- Registers
 has_written_to_t,
 t8,
 device_in_result,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_return_output,
 device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_return_output,
 result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_return_output,
 t8_MUX_uxn_opcodes_h_l403_c2_b756_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output,
 device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output,
 t8_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output,
 sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l424_c9_dde0_return_output,
 MUX_uxn_opcodes_h_l424_c9_6298_return_output,
 UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8f5f_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_return_output,
 device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l426_c37_889a_return_output,
 device_in_uxn_opcodes_h_l426_c23_b350_return_output,
 UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2186_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : device_in_result_t;
 variable VAR_device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6_uxn_opcodes_h_l403_c2_b756_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l414_c3_85b8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l408_c3_43e7 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l403_c2_b756_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l403_c2_b756_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l403_c2_b756_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l403_c2_b756_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_cond : unsigned(0 downto 0);
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l423_c3_ff58 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l419_c7_e8d9_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l424_c9_6298_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_dde0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_dde0_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_dde0_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l424_c9_6298_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l424_c9_6298_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l424_c9_6298_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d_uxn_opcodes_h_l425_c8_32ce_return_output : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8f5f_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8f5f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_cond : unsigned(0 downto 0);
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_iftrue : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_iffalse : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_cond : unsigned(0 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_b350_device_address : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_b350_phase : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_b350_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_889a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_889a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_889a_return_output : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_b350_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_b350_return_output : device_in_result_t;
 variable VAR_CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d_uxn_opcodes_h_l427_c32_8b83_return_output : unsigned(7 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2186_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2186_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l431_c5_8423 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d_uxn_opcodes_h_l432_c23_68aa_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l403_l429_l419_l425_DUPLICATE_724f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l403_l419_l425_DUPLICATE_1bbe_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l429_l419_l425_DUPLICATE_d713_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l419_l425_DUPLICATE_cf01_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l429_l419_l425_DUPLICATE_cee7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8fbf_uxn_opcodes_h_l441_l397_DUPLICATE_845d_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_has_written_to_t : unsigned(0 downto 0);
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_device_in_result : device_in_result_t;
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_has_written_to_t := has_written_to_t;
  REG_VAR_t8 := t8;
  REG_VAR_device_in_result := device_in_result;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_dde0_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l431_c5_8423 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l431_c5_8423;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_iftrue := to_unsigned(0, 1);
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue := to_unsigned(1, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l423_c3_ff58 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse := VAR_result_sp_relative_shift_uxn_opcodes_h_l423_c3_ff58;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_iftrue := to_unsigned(0, 1);
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_iftrue := to_unsigned(0, 1);
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l408_c3_43e7 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l408_c3_43e7;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l414_c3_85b8 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l414_c3_85b8;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_889a_right := to_unsigned(2, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_right := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_device_ram_read := previous_device_ram_read;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse := VAR_CLOCK_ENABLE;
     VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue := device_in_result;
     VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_iffalse := device_in_result;
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2186_expr := has_written_to_t;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue := has_written_to_t;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_iftrue := has_written_to_t;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse := has_written_to_t;
     VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_dde0_left := VAR_phase;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_889a_left := VAR_phase;
     VAR_device_in_uxn_opcodes_h_l426_c23_b350_previous_device_ram_read := VAR_previous_device_ram_read;
     VAR_MUX_uxn_opcodes_h_l424_c9_6298_iftrue := VAR_previous_stack_read;
     VAR_MUX_uxn_opcodes_h_l424_c9_6298_iffalse := t8;
     VAR_t8_MUX_uxn_opcodes_h_l403_c2_b756_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue := t8;
     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l403_c2_b756] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l403_c2_b756_return_output := result.is_vram_write;

     -- UNARY_OP_NOT[uxn_opcodes_h_l429_c9_2186] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2186_expr <= VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2186_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2186_return_output := UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2186_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l403_l419_l425_DUPLICATE_1bbe LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l403_l419_l425_DUPLICATE_1bbe_return_output := result.device_ram_address;

     -- device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6[uxn_opcodes_h_l403_c2_b756] LATENCY=0
     VAR_device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6_uxn_opcodes_h_l403_c2_b756_return_output := CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6(
     device_in_result,
     to_unsigned(0, 1));

     -- BIN_OP_MINUS[uxn_opcodes_h_l426_c37_889a] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l426_c37_889a_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_889a_left;
     BIN_OP_MINUS_uxn_opcodes_h_l426_c37_889a_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_889a_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_889a_return_output := BIN_OP_MINUS_uxn_opcodes_h_l426_c37_889a_return_output;

     -- CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d[uxn_opcodes_h_l432_c23_68aa] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d_uxn_opcodes_h_l432_c23_68aa_return_output := device_in_result.dei_value;

     -- result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d[uxn_opcodes_h_l403_c2_b756] LATENCY=0
     VAR_result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l403_c2_b756_return_output := result.is_device_ram_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l403_c2_b756] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l403_c2_b756_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d[uxn_opcodes_h_l425_c8_32ce] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d_uxn_opcodes_h_l425_c8_32ce_return_output := device_in_result.is_dei_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l403_c6_2848] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_left;
     BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_return_output := BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l419_c11_29ea] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_left;
     BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_return_output := BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l403_c2_b756] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l403_c2_b756_return_output := result.is_ram_write;

     -- sp_relative_shift[uxn_opcodes_h_l420_c30_0a72] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_ins;
     sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_x <= VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_x;
     sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_y <= VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_return_output := sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l424_c9_dde0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l424_c9_dde0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_dde0_left;
     BIN_OP_EQ_uxn_opcodes_h_l424_c9_dde0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_dde0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_dde0_return_output := BIN_OP_EQ_uxn_opcodes_h_l424_c9_dde0_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l429_l419_l425_DUPLICATE_d713 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l429_l419_l425_DUPLICATE_d713_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l429_l419_l425_DUPLICATE_cee7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l429_l419_l425_DUPLICATE_cee7_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l419_l425_DUPLICATE_cf01 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l419_l425_DUPLICATE_cf01_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l403_l429_l419_l425_DUPLICATE_724f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l403_l429_l419_l425_DUPLICATE_724f_return_output := result.u8_value;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l403_c2_b756] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l403_c2_b756_return_output := result.is_stack_index_flipped;

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l403_c2_b756_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_2848_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l419_c7_e8d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_29ea_return_output;
     VAR_MUX_uxn_opcodes_h_l424_c9_6298_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_dde0_return_output;
     VAR_device_in_uxn_opcodes_h_l426_c23_b350_phase := VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_889a_return_output;
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8f5f_expr := VAR_CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d_uxn_opcodes_h_l425_c8_32ce_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l429_l419_l425_DUPLICATE_cee7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l429_l419_l425_DUPLICATE_cee7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l429_l419_l425_DUPLICATE_cee7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l419_l425_DUPLICATE_cf01_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l419_l425_DUPLICATE_cf01_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l429_l419_l425_DUPLICATE_d713_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l429_l419_l425_DUPLICATE_d713_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l429_l419_l425_DUPLICATE_d713_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue := VAR_CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d_uxn_opcodes_h_l432_c23_68aa_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l403_l419_l425_DUPLICATE_1bbe_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l403_l419_l425_DUPLICATE_1bbe_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l403_l419_l425_DUPLICATE_1bbe_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l403_l429_l419_l425_DUPLICATE_724f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l403_l429_l419_l425_DUPLICATE_724f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l403_l429_l419_l425_DUPLICATE_724f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l403_l429_l419_l425_DUPLICATE_724f_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2186_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2186_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2186_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2186_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2186_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_iftrue := VAR_device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6_uxn_opcodes_h_l403_c2_b756_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_iffalse := VAR_result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l403_c2_b756_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l403_c2_b756_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l403_c2_b756_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l403_c2_b756_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l403_c2_b756_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_0a72_return_output;
     -- result_is_device_ram_write_MUX[uxn_opcodes_h_l403_c2_b756] LATENCY=0
     -- Inputs
     result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_cond <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_cond;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_iftrue <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_iftrue;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_iffalse <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_iffalse;
     -- Outputs
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output := result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l403_c2_b756] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l403_c2_b756] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l429_c4_e1db] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l403_c2_b756] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_return_output;

     -- UNARY_OP_NOT[uxn_opcodes_h_l425_c8_8f5f] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8f5f_expr <= VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8f5f_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8f5f_return_output := UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8f5f_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l419_c7_e8d9] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l419_c7_e8d9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l429_c4_e1db] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l429_c4_e1db] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_cond;
     result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_return_output := result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l403_c2_b756] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l429_c4_e1db] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_return_output := has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l429_c4_e1db] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_return_output;

     -- MUX[uxn_opcodes_h_l424_c9_6298] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l424_c9_6298_cond <= VAR_MUX_uxn_opcodes_h_l424_c9_6298_cond;
     MUX_uxn_opcodes_h_l424_c9_6298_iftrue <= VAR_MUX_uxn_opcodes_h_l424_c9_6298_iftrue;
     MUX_uxn_opcodes_h_l424_c9_6298_iffalse <= VAR_MUX_uxn_opcodes_h_l424_c9_6298_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l424_c9_6298_return_output := MUX_uxn_opcodes_h_l424_c9_6298_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output;
     VAR_device_in_uxn_opcodes_h_l426_c23_b350_device_address := VAR_MUX_uxn_opcodes_h_l424_c9_6298_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse := VAR_MUX_uxn_opcodes_h_l424_c9_6298_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8f5f_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8f5f_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8f5f_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8f5f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8f5f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8f5f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8f5f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_8f5f_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_iffalse := VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_e1db_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_e1db_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_e1db_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_e1db_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_e1db_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l403_c2_b756] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l422_c1_340c] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l425_c3_8930] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_return_output := has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l425_c3_8930] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_return_output;

     -- t8_MUX[uxn_opcodes_h_l419_c7_e8d9] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l419_c7_e8d9_cond <= VAR_t8_MUX_uxn_opcodes_h_l419_c7_e8d9_cond;
     t8_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue;
     t8_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output := t8_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l425_c3_8930] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l425_c3_8930] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l425_c3_8930] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_cond;
     result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_return_output := result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_return_output;

     -- Submodule level 3
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_340c_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse := VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_8930_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_8930_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_8930_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_8930_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_8930_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l403_c2_b756_iffalse := VAR_t8_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l419_c7_e8d9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output := result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l425_c1_46c8] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l419_c7_e8d9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l419_c7_e8d9] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output := has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l419_c7_e8d9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l419_c7_e8d9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output;

     -- t8_MUX[uxn_opcodes_h_l403_c2_b756] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l403_c2_b756_cond <= VAR_t8_MUX_uxn_opcodes_h_l403_c2_b756_cond;
     t8_MUX_uxn_opcodes_h_l403_c2_b756_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l403_c2_b756_iftrue;
     t8_MUX_uxn_opcodes_h_l403_c2_b756_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l403_c2_b756_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l403_c2_b756_return_output := t8_MUX_uxn_opcodes_h_l403_c2_b756_return_output;

     -- Submodule level 4
     VAR_device_in_uxn_opcodes_h_l426_c23_b350_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_46c8_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_iffalse := VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l403_c2_b756_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l403_c2_b756] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l403_c2_b756] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l403_c2_b756] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l403_c2_b756] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_return_output := has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_return_output;

     -- device_in[uxn_opcodes_h_l426_c23_b350] LATENCY=0
     -- Clock enable
     device_in_uxn_opcodes_h_l426_c23_b350_CLOCK_ENABLE <= VAR_device_in_uxn_opcodes_h_l426_c23_b350_CLOCK_ENABLE;
     -- Inputs
     device_in_uxn_opcodes_h_l426_c23_b350_device_address <= VAR_device_in_uxn_opcodes_h_l426_c23_b350_device_address;
     device_in_uxn_opcodes_h_l426_c23_b350_phase <= VAR_device_in_uxn_opcodes_h_l426_c23_b350_phase;
     device_in_uxn_opcodes_h_l426_c23_b350_previous_device_ram_read <= VAR_device_in_uxn_opcodes_h_l426_c23_b350_previous_device_ram_read;
     -- Outputs
     VAR_device_in_uxn_opcodes_h_l426_c23_b350_return_output := device_in_uxn_opcodes_h_l426_c23_b350_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l403_c2_b756] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_cond;
     result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_return_output := result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_return_output;

     -- Submodule level 5
     VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_iftrue := VAR_device_in_uxn_opcodes_h_l426_c23_b350_return_output;
     REG_VAR_has_written_to_t := VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_b756_return_output;
     -- device_in_result_MUX[uxn_opcodes_h_l425_c3_8930] LATENCY=0
     -- Inputs
     device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_cond <= VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_cond;
     device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_iftrue <= VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_iftrue;
     device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_iffalse <= VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_iffalse;
     -- Outputs
     VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_return_output := device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_return_output;

     -- CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d[uxn_opcodes_h_l427_c32_8b83] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d_uxn_opcodes_h_l427_c32_8b83_return_output := VAR_device_in_uxn_opcodes_h_l426_c23_b350_return_output.device_ram_address;

     -- Submodule level 6
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_iftrue := VAR_CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d_uxn_opcodes_h_l427_c32_8b83_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse := VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_8930_return_output;
     -- result_device_ram_address_MUX[uxn_opcodes_h_l425_c3_8930] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_return_output;

     -- device_in_result_MUX[uxn_opcodes_h_l419_c7_e8d9] LATENCY=0
     -- Inputs
     device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_cond <= VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_cond;
     device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue <= VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue;
     device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse <= VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse;
     -- Outputs
     VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output := device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output;

     -- Submodule level 7
     VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_iffalse := VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_8930_return_output;
     -- result_device_ram_address_MUX[uxn_opcodes_h_l419_c7_e8d9] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output;

     -- device_in_result_MUX[uxn_opcodes_h_l403_c2_b756] LATENCY=0
     -- Inputs
     device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_cond <= VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_cond;
     device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_iftrue <= VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_iftrue;
     device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_iffalse <= VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_iffalse;
     -- Outputs
     VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_return_output := device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_return_output;

     -- Submodule level 8
     REG_VAR_device_in_result := VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_b756_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_e8d9_return_output;
     -- result_device_ram_address_MUX[uxn_opcodes_h_l403_c2_b756] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_return_output;

     -- Submodule level 9
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8fbf_uxn_opcodes_h_l441_l397_DUPLICATE_845d LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8fbf_uxn_opcodes_h_l441_l397_DUPLICATE_845d_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8fbf(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_b756_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_b756_return_output,
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_b756_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_b756_return_output,
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_b756_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_b756_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_b756_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_b756_return_output);

     -- Submodule level 10
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8fbf_uxn_opcodes_h_l441_l397_DUPLICATE_845d_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8fbf_uxn_opcodes_h_l441_l397_DUPLICATE_845d_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_has_written_to_t <= REG_VAR_has_written_to_t;
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_device_in_result <= REG_VAR_device_in_result;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     has_written_to_t <= REG_COMB_has_written_to_t;
     t8 <= REG_COMB_t8;
     device_in_result <= REG_COMB_device_in_result;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
