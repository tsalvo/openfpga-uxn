-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 50
entity ldr_0CLK_b128164d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldr_0CLK_b128164d;
architecture arch of ldr_0CLK_b128164d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1416_c6_ba57]
signal BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1416_c2_9367]
signal tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1416_c2_9367]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1416_c2_9367]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1416_c2_9367]
signal result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1416_c2_9367]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1416_c2_9367]
signal result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1416_c2_9367]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1416_c2_9367]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1416_c2_9367]
signal t8_MUX_uxn_opcodes_h_l1416_c2_9367_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1416_c2_9367_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1423_c11_b00a]
signal BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1423_c7_34c2]
signal tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1423_c7_34c2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1423_c7_34c2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1423_c7_34c2]
signal result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1423_c7_34c2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1423_c7_34c2]
signal result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1423_c7_34c2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1423_c7_34c2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1423_c7_34c2]
signal t8_MUX_uxn_opcodes_h_l1423_c7_34c2_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1426_c11_0443]
signal BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1426_c7_7b3b]
signal tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1426_c7_7b3b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1426_c7_7b3b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1426_c7_7b3b]
signal result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1426_c7_7b3b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1426_c7_7b3b]
signal result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1426_c7_7b3b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1426_c7_7b3b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1426_c7_7b3b]
signal t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1429_c30_3b62]
signal sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_return_output : signed(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1430_c22_a157]
signal BIN_OP_PLUS_uxn_opcodes_h_l1430_c22_a157_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1430_c22_a157_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1430_c22_a157_return_output : signed(17 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1432_c11_2bd0]
signal BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1432_c7_8e0a]
signal tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1432_c7_8e0a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1432_c7_8e0a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1432_c7_8e0a]
signal result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1432_c7_8e0a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1432_c7_8e0a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1435_c11_7d4c]
signal BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1435_c7_9560]
signal tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1435_c7_9560]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1435_c7_9560]
signal result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1435_c7_9560]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1435_c7_9560]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1441_c11_20be]
signal BIN_OP_EQ_uxn_opcodes_h_l1441_c11_20be_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1441_c11_20be_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1441_c11_20be_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1441_c7_c319]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1441_c7_c319]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_return_output : unsigned(0 downto 0);

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_44b7( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_stack_write := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57
BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_left,
BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_right,
BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1416_c2_9367
tmp8_MUX_uxn_opcodes_h_l1416_c2_9367 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_cond,
tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue,
tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse,
tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367
result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367
result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_cond,
result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367
result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367
result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_cond,
result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367
result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367
result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_return_output);

-- t8_MUX_uxn_opcodes_h_l1416_c2_9367
t8_MUX_uxn_opcodes_h_l1416_c2_9367 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1416_c2_9367_cond,
t8_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue,
t8_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse,
t8_MUX_uxn_opcodes_h_l1416_c2_9367_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a
BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_left,
BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_right,
BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2
tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_cond,
tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue,
tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse,
tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2
result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2
result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_cond,
result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2
result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2
result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_cond,
result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2
result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2
result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output);

-- t8_MUX_uxn_opcodes_h_l1423_c7_34c2
t8_MUX_uxn_opcodes_h_l1423_c7_34c2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1423_c7_34c2_cond,
t8_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue,
t8_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse,
t8_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443
BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_left,
BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_right,
BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b
tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond,
tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue,
tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse,
tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b
result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b
result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond,
result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b
result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b
result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b
result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output);

-- t8_MUX_uxn_opcodes_h_l1426_c7_7b3b
t8_MUX_uxn_opcodes_h_l1426_c7_7b3b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond,
t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue,
t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse,
t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62
sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_ins,
sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_x,
sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_y,
sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1430_c22_a157
BIN_OP_PLUS_uxn_opcodes_h_l1430_c22_a157 : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1430_c22_a157_left,
BIN_OP_PLUS_uxn_opcodes_h_l1430_c22_a157_right,
BIN_OP_PLUS_uxn_opcodes_h_l1430_c22_a157_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0
BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0_left,
BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0_right,
BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a
tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond,
tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue,
tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse,
tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a
result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a
result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a
result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond,
result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a
result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c
BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c_left,
BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c_right,
BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1435_c7_9560
tmp8_MUX_uxn_opcodes_h_l1435_c7_9560 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_cond,
tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue,
tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse,
tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560
result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560
result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_cond,
result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560
result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1441_c11_20be
BIN_OP_EQ_uxn_opcodes_h_l1441_c11_20be : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1441_c11_20be_left,
BIN_OP_EQ_uxn_opcodes_h_l1441_c11_20be_right,
BIN_OP_EQ_uxn_opcodes_h_l1441_c11_20be_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319
result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319
result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_return_output,
 tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_return_output,
 t8_MUX_uxn_opcodes_h_l1416_c2_9367_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_return_output,
 tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output,
 t8_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_return_output,
 tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output,
 t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output,
 sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1430_c22_a157_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0_return_output,
 tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c_return_output,
 tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1441_c11_20be_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1420_c3_d558 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1416_c2_9367_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1416_c2_9367_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1424_c3_c0ea : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1423_c7_34c2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l1430_c3_a703 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1430_c22_a157_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l1430_c27_3433_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1430_c22_a157_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1430_c22_a157_return_output : signed(17 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1438_c3_96f3 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_20be_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_20be_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_20be_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1423_l1416_l1432_DUPLICATE_dd14_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1423_l1426_l1416_DUPLICATE_3f0c_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1423_l1416_l1435_l1432_l1426_DUPLICATE_f5b6_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1423_l1426_l1416_DUPLICATE_54ce_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1423_l1416_l1432_l1441_l1426_DUPLICATE_0c7c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1423_l1435_l1432_l1441_l1426_DUPLICATE_3544_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1435_l1426_l1432_DUPLICATE_2185_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_44b7_uxn_opcodes_h_l1412_l1446_DUPLICATE_5c07_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1438_c3_96f3 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1438_c3_96f3;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1420_c3_d558 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1420_c3_d558;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_20be_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1424_c3_c0ea := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1424_c3_c0ea;
     VAR_sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_ins := VAR_ins;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1430_c22_a157_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_20be_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse := tmp8;
     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1435_l1426_l1432_DUPLICATE_2185 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1435_l1426_l1432_DUPLICATE_2185_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1423_l1426_l1416_DUPLICATE_3f0c LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1423_l1426_l1416_DUPLICATE_3f0c_return_output := result.u16_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1432_c11_2bd0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0_left;
     BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0_return_output := BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1423_l1416_l1435_l1432_l1426_DUPLICATE_f5b6 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1423_l1416_l1435_l1432_l1426_DUPLICATE_f5b6_return_output := result.u8_value;

     -- CAST_TO_int8_t[uxn_opcodes_h_l1430_c27_3433] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l1430_c27_3433_return_output := CAST_TO_int8_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l1435_c11_7d4c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1423_l1416_l1432_DUPLICATE_dd14 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1423_l1416_l1432_DUPLICATE_dd14_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1441_c11_20be] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1441_c11_20be_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_20be_left;
     BIN_OP_EQ_uxn_opcodes_h_l1441_c11_20be_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_20be_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_20be_return_output := BIN_OP_EQ_uxn_opcodes_h_l1441_c11_20be_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1423_l1426_l1416_DUPLICATE_54ce LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1423_l1426_l1416_DUPLICATE_54ce_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1416_c6_ba57] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_left;
     BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_return_output := BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1426_c11_0443] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_left;
     BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_return_output := BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1429_c30_3b62] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_ins;
     sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_x;
     sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_return_output := sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1423_c11_b00a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1423_l1435_l1432_l1441_l1426_DUPLICATE_3544 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1423_l1435_l1432_l1441_l1426_DUPLICATE_3544_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1423_l1416_l1432_l1441_l1426_DUPLICATE_0c7c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1423_l1416_l1432_l1441_l1426_DUPLICATE_0c7c_return_output := result.is_stack_write;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1416_c2_9367_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c6_ba57_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1423_c7_34c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1423_c11_b00a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1426_c11_0443_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1432_c11_2bd0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1435_c11_7d4c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_20be_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1441_c11_20be_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1430_c22_a157_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l1430_c27_3433_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1423_l1426_l1416_DUPLICATE_54ce_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1423_l1426_l1416_DUPLICATE_54ce_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1423_l1426_l1416_DUPLICATE_54ce_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1423_l1426_l1416_DUPLICATE_3f0c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1423_l1426_l1416_DUPLICATE_3f0c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1423_l1426_l1416_DUPLICATE_3f0c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1423_l1435_l1432_l1441_l1426_DUPLICATE_3544_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1423_l1435_l1432_l1441_l1426_DUPLICATE_3544_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1423_l1435_l1432_l1441_l1426_DUPLICATE_3544_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1423_l1435_l1432_l1441_l1426_DUPLICATE_3544_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1423_l1435_l1432_l1441_l1426_DUPLICATE_3544_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1423_l1416_l1432_DUPLICATE_dd14_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1423_l1416_l1432_DUPLICATE_dd14_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1423_l1416_l1432_DUPLICATE_dd14_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1423_l1416_l1432_l1441_l1426_DUPLICATE_0c7c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1423_l1416_l1432_l1441_l1426_DUPLICATE_0c7c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1423_l1416_l1432_l1441_l1426_DUPLICATE_0c7c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1423_l1416_l1432_l1441_l1426_DUPLICATE_0c7c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1423_l1416_l1432_l1441_l1426_DUPLICATE_0c7c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1435_l1426_l1432_DUPLICATE_2185_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1435_l1426_l1432_DUPLICATE_2185_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1435_l1426_l1432_DUPLICATE_2185_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1423_l1416_l1435_l1432_l1426_DUPLICATE_f5b6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1423_l1416_l1435_l1432_l1426_DUPLICATE_f5b6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1423_l1416_l1435_l1432_l1426_DUPLICATE_f5b6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1423_l1416_l1435_l1432_l1426_DUPLICATE_f5b6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1423_l1416_l1435_l1432_l1426_DUPLICATE_f5b6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1429_c30_3b62_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l1435_c7_9560] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_cond;
     tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_return_output := tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1426_c7_7b3b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1432_c7_8e0a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1430_c22_a157] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1430_c22_a157_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1430_c22_a157_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1430_c22_a157_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1430_c22_a157_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1430_c22_a157_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1430_c22_a157_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1441_c7_c319] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_return_output;

     -- t8_MUX[uxn_opcodes_h_l1426_c7_7b3b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond <= VAR_t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond;
     t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue;
     t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output := t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1441_c7_c319] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1435_c7_9560] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1435_c7_9560] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_return_output := result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_return_output;

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l1430_c3_a703 := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1430_c22_a157_return_output)),16);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1441_c7_c319_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1441_c7_c319_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1435_c7_9560_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1435_c7_9560_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1435_c7_9560_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue := VAR_result_u16_value_uxn_opcodes_h_l1430_c3_a703;
     -- tmp8_MUX[uxn_opcodes_h_l1432_c7_8e0a] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond;
     tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output := tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1432_c7_8e0a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output := result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1423_c7_34c2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1435_c7_9560] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1435_c7_9560] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_return_output;

     -- t8_MUX[uxn_opcodes_h_l1423_c7_34c2] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1423_c7_34c2_cond <= VAR_t8_MUX_uxn_opcodes_h_l1423_c7_34c2_cond;
     t8_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue;
     t8_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output := t8_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1426_c7_7b3b] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output := result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1432_c7_8e0a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1426_c7_7b3b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1435_c7_9560_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1435_c7_9560_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output;
     -- t8_MUX[uxn_opcodes_h_l1416_c2_9367] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1416_c2_9367_cond <= VAR_t8_MUX_uxn_opcodes_h_l1416_c2_9367_cond;
     t8_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue;
     t8_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1416_c2_9367_return_output := t8_MUX_uxn_opcodes_h_l1416_c2_9367_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1416_c2_9367] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1426_c7_7b3b] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond;
     tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output := tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1426_c7_7b3b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1423_c7_34c2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1432_c7_8e0a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1423_c7_34c2] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output := result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1426_c7_7b3b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1432_c7_8e0a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1432_c7_8e0a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1416_c2_9367_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l1423_c7_34c2] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_cond;
     tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output := tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1426_c7_7b3b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1416_c2_9367] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1423_c7_34c2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1426_c7_7b3b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1423_c7_34c2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output := result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1416_c2_9367] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_return_output := result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1426_c7_7b3b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l1416_c2_9367] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_cond;
     tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_return_output := tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1416_c2_9367] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1423_c7_34c2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1416_c2_9367] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_return_output := result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1423_c7_34c2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1423_c7_34c2_return_output;
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1416_c2_9367_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1416_c2_9367] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1416_c2_9367] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_44b7_uxn_opcodes_h_l1412_l1446_DUPLICATE_5c07 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_44b7_uxn_opcodes_h_l1412_l1446_DUPLICATE_5c07_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_44b7(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c2_9367_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1416_c2_9367_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1416_c2_9367_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1416_c2_9367_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1416_c2_9367_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c2_9367_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1416_c2_9367_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_44b7_uxn_opcodes_h_l1412_l1446_DUPLICATE_5c07_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_44b7_uxn_opcodes_h_l1412_l1446_DUPLICATE_5c07_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
