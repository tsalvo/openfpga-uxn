-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 57
entity jsr2_0CLK_609876da is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jsr2_0CLK_609876da;
architecture arch of jsr2_0CLK_609876da is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l773_c6_65c0]
signal BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l773_c2_b814]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l773_c2_b814]
signal result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l773_c2_b814]
signal result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l773_c2_b814]
signal result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l773_c2_b814]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l773_c2_b814]
signal result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l773_c2_b814]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l773_c2_b814]
signal result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l773_c2_b814]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l773_c2_b814]
signal result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l773_c2_b814]
signal t16_MUX_uxn_opcodes_h_l773_c2_b814_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l773_c2_b814_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l773_c2_b814_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l773_c2_b814_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l786_c11_5d1f]
signal BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l786_c7_d4c9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l786_c7_d4c9]
signal result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l786_c7_d4c9]
signal result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output : unsigned(15 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l786_c7_d4c9]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l786_c7_d4c9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l786_c7_d4c9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l786_c7_d4c9]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l786_c7_d4c9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l786_c7_d4c9]
signal t16_MUX_uxn_opcodes_h_l786_c7_d4c9_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l789_c11_89b2]
signal BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l789_c7_4356]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l789_c7_4356]
signal result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l789_c7_4356]
signal result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_return_output : unsigned(15 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l789_c7_4356]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l789_c7_4356]
signal result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l789_c7_4356]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l789_c7_4356]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l789_c7_4356]
signal result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l789_c7_4356]
signal t16_MUX_uxn_opcodes_h_l789_c7_4356_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l789_c7_4356_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l789_c7_4356_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l789_c7_4356_return_output : unsigned(15 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l791_c3_8fad]
signal CONST_SL_8_uxn_opcodes_h_l791_c3_8fad_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l791_c3_8fad_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l792_c30_24b6]
signal sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l794_c11_54c2]
signal BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l794_c7_52e3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l794_c7_52e3]
signal result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l794_c7_52e3]
signal result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_return_output : unsigned(15 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l794_c7_52e3]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l794_c7_52e3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l794_c7_52e3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l794_c7_52e3]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l794_c7_52e3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l794_c7_52e3]
signal t16_MUX_uxn_opcodes_h_l794_c7_52e3_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l794_c7_52e3_return_output : unsigned(15 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l795_c3_6d5d]
signal BIN_OP_OR_uxn_opcodes_h_l795_c3_6d5d_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l795_c3_6d5d_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l795_c3_6d5d_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l802_c11_fe8d]
signal BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l802_c7_a1f7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l802_c7_a1f7]
signal result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l802_c7_a1f7]
signal result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l802_c7_a1f7]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l802_c7_a1f7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l802_c7_a1f7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output : unsigned(0 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l805_c31_a93c]
signal CONST_SR_8_uxn_opcodes_h_l805_c31_a93c_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l805_c31_a93c_return_output : unsigned(15 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_e393( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_ram_write := ref_toks_4;
      base.is_stack_index_flipped := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_vram_write := ref_toks_8;
      base.is_pc_updated := ref_toks_9;
      base.is_opc_done := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0
BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_left,
BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_right,
BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814
result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_cond,
result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814
result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_cond,
result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814
result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814
result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814
result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814
result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814
result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814
result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_return_output);

-- t16_MUX_uxn_opcodes_h_l773_c2_b814
t16_MUX_uxn_opcodes_h_l773_c2_b814 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l773_c2_b814_cond,
t16_MUX_uxn_opcodes_h_l773_c2_b814_iftrue,
t16_MUX_uxn_opcodes_h_l773_c2_b814_iffalse,
t16_MUX_uxn_opcodes_h_l773_c2_b814_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f
BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_left,
BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_right,
BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9
result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_cond,
result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9
result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_cond,
result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9
result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9
result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9
result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9
result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output);

-- t16_MUX_uxn_opcodes_h_l786_c7_d4c9
t16_MUX_uxn_opcodes_h_l786_c7_d4c9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l786_c7_d4c9_cond,
t16_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue,
t16_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse,
t16_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2
BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_left,
BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_right,
BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356
result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_cond,
result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356
result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_cond,
result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356
result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356
result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356
result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356
result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_return_output);

-- t16_MUX_uxn_opcodes_h_l789_c7_4356
t16_MUX_uxn_opcodes_h_l789_c7_4356 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l789_c7_4356_cond,
t16_MUX_uxn_opcodes_h_l789_c7_4356_iftrue,
t16_MUX_uxn_opcodes_h_l789_c7_4356_iffalse,
t16_MUX_uxn_opcodes_h_l789_c7_4356_return_output);

-- CONST_SL_8_uxn_opcodes_h_l791_c3_8fad
CONST_SL_8_uxn_opcodes_h_l791_c3_8fad : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l791_c3_8fad_x,
CONST_SL_8_uxn_opcodes_h_l791_c3_8fad_return_output);

-- sp_relative_shift_uxn_opcodes_h_l792_c30_24b6
sp_relative_shift_uxn_opcodes_h_l792_c30_24b6 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_ins,
sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_x,
sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_y,
sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2
BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_left,
BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_right,
BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3
result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_cond,
result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3
result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_cond,
result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3
result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3
result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3
result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3
result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_return_output);

-- t16_MUX_uxn_opcodes_h_l794_c7_52e3
t16_MUX_uxn_opcodes_h_l794_c7_52e3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l794_c7_52e3_cond,
t16_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue,
t16_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse,
t16_MUX_uxn_opcodes_h_l794_c7_52e3_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l795_c3_6d5d
BIN_OP_OR_uxn_opcodes_h_l795_c3_6d5d : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l795_c3_6d5d_left,
BIN_OP_OR_uxn_opcodes_h_l795_c3_6d5d_right,
BIN_OP_OR_uxn_opcodes_h_l795_c3_6d5d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d
BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d_left,
BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d_right,
BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7
result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_cond,
result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7
result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_cond,
result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7
result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7
result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7
result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output);

-- CONST_SR_8_uxn_opcodes_h_l805_c31_a93c
CONST_SR_8_uxn_opcodes_h_l805_c31_a93c : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l805_c31_a93c_x,
CONST_SR_8_uxn_opcodes_h_l805_c31_a93c_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 -- Registers
 t16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_return_output,
 t16_MUX_uxn_opcodes_h_l773_c2_b814_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output,
 t16_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_return_output,
 t16_MUX_uxn_opcodes_h_l789_c7_4356_return_output,
 CONST_SL_8_uxn_opcodes_h_l791_c3_8fad_return_output,
 sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_return_output,
 t16_MUX_uxn_opcodes_h_l794_c7_52e3_return_output,
 BIN_OP_OR_uxn_opcodes_h_l795_c3_6d5d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output,
 CONST_SR_8_uxn_opcodes_h_l805_c31_a93c_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l783_c3_7af7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l773_c2_b814_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l778_c3_40c0 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l773_c2_b814_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l773_c2_b814_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l773_c2_b814_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l773_c2_b814_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l773_c2_b814_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l787_c3_bc70 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l789_c7_4356_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l786_c7_d4c9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l789_c7_4356_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l789_c7_4356_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l794_c7_52e3_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l789_c7_4356_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l791_c3_8fad_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l791_c3_8fad_x : unsigned(15 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l799_c3_f1d7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l797_c3_e730 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l794_c7_52e3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l795_c3_6d5d_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l795_c3_6d5d_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l795_c3_6d5d_return_output : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l800_c21_8be2_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l804_c3_f832 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l803_c3_9a29 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l805_c31_a93c_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l805_c31_a93c_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l805_c21_a5b1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l789_l773_l786_l802_DUPLICATE_14e6_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l789_l773_l802_l794_l786_DUPLICATE_511f_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l794_l789_l786_DUPLICATE_7d77_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l794_l789_l786_DUPLICATE_c359_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l786_l802_DUPLICATE_be2e_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l794_l789_l786_l802_DUPLICATE_802d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l794_l789_l786_l802_DUPLICATE_3022_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l790_l795_DUPLICATE_3fe0_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l789_l802_DUPLICATE_13b8_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e393_uxn_opcodes_h_l811_l769_DUPLICATE_9d83_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_y := resize(to_signed(-2, 3), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l804_c3_f832 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l804_c3_f832;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_right := to_unsigned(2, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l803_c3_9a29 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l803_c3_9a29;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_right := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l797_c3_e730 := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l797_c3_e730;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l787_c3_bc70 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l787_c3_bc70;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l799_c3_f1d7 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l799_c3_f1d7;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l778_c3_40c0 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l778_c3_40c0;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l783_c3_7af7 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l783_c3_7af7;
     VAR_sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_right := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_ins := VAR_ins;
     VAR_CONST_SR_8_uxn_opcodes_h_l805_c31_a93c_x := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l795_c3_6d5d_left := t16;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l773_c2_b814_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse := t16;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l794_l789_l786_l802_DUPLICATE_3022 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l794_l789_l786_l802_DUPLICATE_3022_return_output := result.is_opc_done;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l800_c21_8be2] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l800_c21_8be2_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_pc);

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l773_c2_b814] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l773_c2_b814_return_output := result.is_vram_write;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l790_l795_DUPLICATE_3fe0 LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l790_l795_DUPLICATE_3fe0_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l789_l773_l786_l802_DUPLICATE_14e6 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l789_l773_l786_l802_DUPLICATE_14e6_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l773_c6_65c0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_left;
     BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_return_output := BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l789_c11_89b2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_left;
     BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_return_output := BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l794_c11_54c2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_left;
     BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_return_output := BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l792_c30_24b6] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_ins;
     sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_x <= VAR_sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_x;
     sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_y <= VAR_sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_return_output := sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l789_l773_l802_l794_l786_DUPLICATE_511f LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l789_l773_l802_l794_l786_DUPLICATE_511f_return_output := result.u16_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l794_l789_l786_DUPLICATE_c359 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l794_l789_l786_DUPLICATE_c359_return_output := result.is_stack_write;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l773_c2_b814] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l773_c2_b814_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l794_l789_l786_DUPLICATE_7d77 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l794_l789_l786_DUPLICATE_7d77_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l786_l802_DUPLICATE_be2e LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l786_l802_DUPLICATE_be2e_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l786_c11_5d1f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_left;
     BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_return_output := BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l789_l802_DUPLICATE_13b8 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l789_l802_DUPLICATE_13b8_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l794_l789_l786_l802_DUPLICATE_802d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l794_l789_l786_l802_DUPLICATE_802d_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l802_c11_fe8d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d_left;
     BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d_return_output := BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d_return_output;

     -- CONST_SR_8[uxn_opcodes_h_l805_c31_a93c] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l805_c31_a93c_x <= VAR_CONST_SR_8_uxn_opcodes_h_l805_c31_a93c_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l805_c31_a93c_return_output := CONST_SR_8_uxn_opcodes_h_l805_c31_a93c_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l773_c2_b814_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l773_c6_65c0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l786_c7_d4c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l786_c11_5d1f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l789_c7_4356_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l789_c11_89b2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l794_c7_52e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l794_c11_54c2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l802_c11_fe8d_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l795_c3_6d5d_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l790_l795_DUPLICATE_3fe0_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l791_c3_8fad_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l790_l795_DUPLICATE_3fe0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l800_c21_8be2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l786_l802_DUPLICATE_be2e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l786_l802_DUPLICATE_be2e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l789_l773_l802_l794_l786_DUPLICATE_511f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l789_l773_l802_l794_l786_DUPLICATE_511f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l789_l773_l802_l794_l786_DUPLICATE_511f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l789_l773_l802_l794_l786_DUPLICATE_511f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l789_l773_l802_l794_l786_DUPLICATE_511f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l794_l789_l786_l802_DUPLICATE_3022_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l794_l789_l786_l802_DUPLICATE_3022_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l794_l789_l786_l802_DUPLICATE_3022_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l794_l789_l786_l802_DUPLICATE_3022_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l794_l789_l786_l802_DUPLICATE_802d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l794_l789_l786_l802_DUPLICATE_802d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l794_l789_l786_l802_DUPLICATE_802d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l794_l789_l786_l802_DUPLICATE_802d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l794_l789_l786_DUPLICATE_7d77_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l794_l789_l786_DUPLICATE_7d77_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l794_l789_l786_DUPLICATE_7d77_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l794_l789_l786_DUPLICATE_c359_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l794_l789_l786_DUPLICATE_c359_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l794_l789_l786_DUPLICATE_c359_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l789_l802_DUPLICATE_13b8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l789_l802_DUPLICATE_13b8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l789_l773_l786_l802_DUPLICATE_14e6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l789_l773_l786_l802_DUPLICATE_14e6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l789_l773_l786_l802_DUPLICATE_14e6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l789_l773_l786_l802_DUPLICATE_14e6_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l773_c2_b814_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l773_c2_b814_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l792_c30_24b6_return_output;
     -- CONST_SL_8[uxn_opcodes_h_l791_c3_8fad] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l791_c3_8fad_x <= VAR_CONST_SL_8_uxn_opcodes_h_l791_c3_8fad_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l791_c3_8fad_return_output := CONST_SL_8_uxn_opcodes_h_l791_c3_8fad_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l773_c2_b814] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l794_c7_52e3] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l802_c7_a1f7] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l795_c3_6d5d] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l795_c3_6d5d_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l795_c3_6d5d_left;
     BIN_OP_OR_uxn_opcodes_h_l795_c3_6d5d_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l795_c3_6d5d_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l795_c3_6d5d_return_output := BIN_OP_OR_uxn_opcodes_h_l795_c3_6d5d_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l773_c2_b814] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l802_c7_a1f7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l802_c7_a1f7] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_cond;
     result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output := result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l802_c7_a1f7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l802_c7_a1f7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l805_c21_a5b1] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l805_c21_a5b1_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l805_c31_a93c_return_output);

     -- result_is_stack_write_MUX[uxn_opcodes_h_l794_c7_52e3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_return_output;

     -- Submodule level 2
     VAR_t16_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l795_c3_6d5d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l805_c21_a5b1_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l789_c7_4356_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l791_c3_8fad_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l794_c7_52e3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l794_c7_52e3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output;
     -- t16_MUX[uxn_opcodes_h_l794_c7_52e3] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l794_c7_52e3_cond <= VAR_t16_MUX_uxn_opcodes_h_l794_c7_52e3_cond;
     t16_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue;
     t16_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l794_c7_52e3_return_output := t16_MUX_uxn_opcodes_h_l794_c7_52e3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l794_c7_52e3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l789_c7_4356] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l794_c7_52e3] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l794_c7_52e3] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_cond;
     result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_return_output := result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l794_c7_52e3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l789_c7_4356] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l794_c7_52e3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l802_c7_a1f7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output := result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l794_c7_52e3_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l794_c7_52e3_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l789_c7_4356_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l789_c7_4356_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l794_c7_52e3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l794_c7_52e3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l794_c7_52e3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l802_c7_a1f7_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l789_c7_4356_iffalse := VAR_t16_MUX_uxn_opcodes_h_l794_c7_52e3_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l794_c7_52e3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_return_output := result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l786_c7_d4c9] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l789_c7_4356] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l789_c7_4356] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_cond;
     result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_return_output := result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l789_c7_4356] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_return_output;

     -- t16_MUX[uxn_opcodes_h_l789_c7_4356] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l789_c7_4356_cond <= VAR_t16_MUX_uxn_opcodes_h_l789_c7_4356_cond;
     t16_MUX_uxn_opcodes_h_l789_c7_4356_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l789_c7_4356_iftrue;
     t16_MUX_uxn_opcodes_h_l789_c7_4356_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l789_c7_4356_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l789_c7_4356_return_output := t16_MUX_uxn_opcodes_h_l789_c7_4356_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l786_c7_d4c9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l789_c7_4356] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l789_c7_4356] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l789_c7_4356_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l789_c7_4356_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l789_c7_4356_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l789_c7_4356_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l789_c7_4356_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l794_c7_52e3_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse := VAR_t16_MUX_uxn_opcodes_h_l789_c7_4356_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l773_c2_b814] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l786_c7_d4c9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l786_c7_d4c9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l786_c7_d4c9] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l786_c7_d4c9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output;

     -- t16_MUX[uxn_opcodes_h_l786_c7_d4c9] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l786_c7_d4c9_cond <= VAR_t16_MUX_uxn_opcodes_h_l786_c7_d4c9_cond;
     t16_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue;
     t16_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output := t16_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l786_c7_d4c9] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_cond;
     result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output := result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l773_c2_b814] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l789_c7_4356] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_cond;
     result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_return_output := result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l789_c7_4356_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l773_c2_b814_iffalse := VAR_t16_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l773_c2_b814] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l773_c2_b814] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l773_c2_b814] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l773_c2_b814] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l773_c2_b814] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_cond;
     result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_return_output := result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_return_output;

     -- t16_MUX[uxn_opcodes_h_l773_c2_b814] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l773_c2_b814_cond <= VAR_t16_MUX_uxn_opcodes_h_l773_c2_b814_cond;
     t16_MUX_uxn_opcodes_h_l773_c2_b814_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l773_c2_b814_iftrue;
     t16_MUX_uxn_opcodes_h_l773_c2_b814_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l773_c2_b814_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l773_c2_b814_return_output := t16_MUX_uxn_opcodes_h_l773_c2_b814_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l786_c7_d4c9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output := result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output;

     -- Submodule level 6
     VAR_result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l786_c7_d4c9_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l773_c2_b814_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l773_c2_b814] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_cond;
     result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_return_output := result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_e393_uxn_opcodes_h_l811_l769_DUPLICATE_9d83 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e393_uxn_opcodes_h_l811_l769_DUPLICATE_9d83_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_e393(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l773_c2_b814_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l773_c2_b814_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l773_c2_b814_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l773_c2_b814_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l773_c2_b814_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l773_c2_b814_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l773_c2_b814_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l773_c2_b814_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l773_c2_b814_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l773_c2_b814_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e393_uxn_opcodes_h_l811_l769_DUPLICATE_9d83_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e393_uxn_opcodes_h_l811_l769_DUPLICATE_9d83_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
