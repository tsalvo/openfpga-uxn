-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity uxn_top_0CLK_8944ffd5 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 is_visible_pixel : in unsigned(0 downto 0);
 rom_load_valid_byte : in unsigned(0 downto 0);
 rom_load_address : in unsigned(15 downto 0);
 rom_load_value : in unsigned(7 downto 0);
 return_output : out unsigned(15 downto 0));
end uxn_top_0CLK_8944ffd5;
architecture arch of uxn_top_0CLK_8944ffd5 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal boot_check : unsigned(23 downto 0) := to_unsigned(0, 24);
signal uxn_eval_result : unsigned(15 downto 0) := to_unsigned(0, 16);
signal is_booted : unsigned(0 downto 0) := to_unsigned(0, 1);
signal gpu_step_result : gpu_step_result_t := gpu_step_result_t_NULL;
signal cpu_step_result : cpu_step_result_t := cpu_step_result_t_NULL;
signal is_active_fill : unsigned(0 downto 0) := to_unsigned(0, 1);
signal is_ram_write : unsigned(0 downto 0) := to_unsigned(0, 1);
signal u16_addr : unsigned(15 downto 0) := to_unsigned(255, 16);
signal screen_vector : unsigned(15 downto 0) := to_unsigned(0, 16);
signal ram_write_value : unsigned(7 downto 0) := to_unsigned(0, 8);
signal ram_read_value : unsigned(7 downto 0) := to_unsigned(0, 8);
signal device_ram_address : unsigned(7 downto 0) := to_unsigned(0, 8);
signal device_ram_read_value : unsigned(7 downto 0) := to_unsigned(0, 8);
signal is_device_ram_write : unsigned(0 downto 0) := to_unsigned(0, 1);
signal is_vram_write : unsigned(0 downto 0) := to_unsigned(0, 1);
signal vram_write_layer : unsigned(0 downto 0) := to_unsigned(0, 1);
signal vram_value : unsigned(7 downto 0) := to_unsigned(0, 8);
signal REG_COMB_boot_check : unsigned(23 downto 0);
signal REG_COMB_uxn_eval_result : unsigned(15 downto 0);
signal REG_COMB_is_booted : unsigned(0 downto 0);
signal REG_COMB_gpu_step_result : gpu_step_result_t;
signal REG_COMB_cpu_step_result : cpu_step_result_t;
signal REG_COMB_is_active_fill : unsigned(0 downto 0);
signal REG_COMB_is_ram_write : unsigned(0 downto 0);
signal REG_COMB_u16_addr : unsigned(15 downto 0);
signal REG_COMB_screen_vector : unsigned(15 downto 0);
signal REG_COMB_ram_write_value : unsigned(7 downto 0);
signal REG_COMB_ram_read_value : unsigned(7 downto 0);
signal REG_COMB_device_ram_address : unsigned(7 downto 0);
signal REG_COMB_device_ram_read_value : unsigned(7 downto 0);
signal REG_COMB_is_device_ram_write : unsigned(0 downto 0);
signal REG_COMB_is_vram_write : unsigned(0 downto 0);
signal REG_COMB_vram_write_layer : unsigned(0 downto 0);
signal REG_COMB_vram_value : unsigned(7 downto 0);

-- Each function instance gets signals
-- UNARY_OP_NOT[uxn_c_l302_c7_51e8]
signal UNARY_OP_NOT_uxn_c_l302_c7_51e8_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_uxn_c_l302_c7_51e8_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_c_l317_c9_9a0e]
signal FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_return_output : unsigned(0 downto 0);

-- u16_addr_MUX[uxn_c_l302_c2_9cba]
signal u16_addr_MUX_uxn_c_l302_c2_9cba_cond : unsigned(0 downto 0);
signal u16_addr_MUX_uxn_c_l302_c2_9cba_iftrue : unsigned(15 downto 0);
signal u16_addr_MUX_uxn_c_l302_c2_9cba_iffalse : unsigned(15 downto 0);
signal u16_addr_MUX_uxn_c_l302_c2_9cba_return_output : unsigned(15 downto 0);

-- vram_write_layer_MUX[uxn_c_l302_c2_9cba]
signal vram_write_layer_MUX_uxn_c_l302_c2_9cba_cond : unsigned(0 downto 0);
signal vram_write_layer_MUX_uxn_c_l302_c2_9cba_iftrue : unsigned(0 downto 0);
signal vram_write_layer_MUX_uxn_c_l302_c2_9cba_iffalse : unsigned(0 downto 0);
signal vram_write_layer_MUX_uxn_c_l302_c2_9cba_return_output : unsigned(0 downto 0);

-- device_ram_address_MUX[uxn_c_l302_c2_9cba]
signal device_ram_address_MUX_uxn_c_l302_c2_9cba_cond : unsigned(0 downto 0);
signal device_ram_address_MUX_uxn_c_l302_c2_9cba_iftrue : unsigned(7 downto 0);
signal device_ram_address_MUX_uxn_c_l302_c2_9cba_iffalse : unsigned(7 downto 0);
signal device_ram_address_MUX_uxn_c_l302_c2_9cba_return_output : unsigned(7 downto 0);

-- is_device_ram_write_MUX[uxn_c_l302_c2_9cba]
signal is_device_ram_write_MUX_uxn_c_l302_c2_9cba_cond : unsigned(0 downto 0);
signal is_device_ram_write_MUX_uxn_c_l302_c2_9cba_iftrue : unsigned(0 downto 0);
signal is_device_ram_write_MUX_uxn_c_l302_c2_9cba_iffalse : unsigned(0 downto 0);
signal is_device_ram_write_MUX_uxn_c_l302_c2_9cba_return_output : unsigned(0 downto 0);

-- is_ram_write_MUX[uxn_c_l302_c2_9cba]
signal is_ram_write_MUX_uxn_c_l302_c2_9cba_cond : unsigned(0 downto 0);
signal is_ram_write_MUX_uxn_c_l302_c2_9cba_iftrue : unsigned(0 downto 0);
signal is_ram_write_MUX_uxn_c_l302_c2_9cba_iffalse : unsigned(0 downto 0);
signal is_ram_write_MUX_uxn_c_l302_c2_9cba_return_output : unsigned(0 downto 0);

-- is_vram_write_MUX[uxn_c_l302_c2_9cba]
signal is_vram_write_MUX_uxn_c_l302_c2_9cba_cond : unsigned(0 downto 0);
signal is_vram_write_MUX_uxn_c_l302_c2_9cba_iftrue : unsigned(0 downto 0);
signal is_vram_write_MUX_uxn_c_l302_c2_9cba_iffalse : unsigned(0 downto 0);
signal is_vram_write_MUX_uxn_c_l302_c2_9cba_return_output : unsigned(0 downto 0);

-- boot_check_MUX[uxn_c_l302_c2_9cba]
signal boot_check_MUX_uxn_c_l302_c2_9cba_cond : unsigned(0 downto 0);
signal boot_check_MUX_uxn_c_l302_c2_9cba_iftrue : unsigned(23 downto 0);
signal boot_check_MUX_uxn_c_l302_c2_9cba_iffalse : unsigned(23 downto 0);
signal boot_check_MUX_uxn_c_l302_c2_9cba_return_output : unsigned(23 downto 0);

-- vram_value_MUX[uxn_c_l302_c2_9cba]
signal vram_value_MUX_uxn_c_l302_c2_9cba_cond : unsigned(0 downto 0);
signal vram_value_MUX_uxn_c_l302_c2_9cba_iftrue : unsigned(7 downto 0);
signal vram_value_MUX_uxn_c_l302_c2_9cba_iffalse : unsigned(7 downto 0);
signal vram_value_MUX_uxn_c_l302_c2_9cba_return_output : unsigned(7 downto 0);

-- ram_write_value_MUX[uxn_c_l302_c2_9cba]
signal ram_write_value_MUX_uxn_c_l302_c2_9cba_cond : unsigned(0 downto 0);
signal ram_write_value_MUX_uxn_c_l302_c2_9cba_iftrue : unsigned(7 downto 0);
signal ram_write_value_MUX_uxn_c_l302_c2_9cba_iffalse : unsigned(7 downto 0);
signal ram_write_value_MUX_uxn_c_l302_c2_9cba_return_output : unsigned(7 downto 0);

-- cpu_step_result_MUX[uxn_c_l302_c2_9cba]
signal cpu_step_result_MUX_uxn_c_l302_c2_9cba_cond : unsigned(0 downto 0);
signal cpu_step_result_MUX_uxn_c_l302_c2_9cba_iftrue : cpu_step_result_t;
signal cpu_step_result_MUX_uxn_c_l302_c2_9cba_iffalse : cpu_step_result_t;
signal cpu_step_result_MUX_uxn_c_l302_c2_9cba_return_output : cpu_step_result_t;

-- is_booted_MUX[uxn_c_l302_c2_9cba]
signal is_booted_MUX_uxn_c_l302_c2_9cba_cond : unsigned(0 downto 0);
signal is_booted_MUX_uxn_c_l302_c2_9cba_iftrue : unsigned(0 downto 0);
signal is_booted_MUX_uxn_c_l302_c2_9cba_iffalse : unsigned(0 downto 0);
signal is_booted_MUX_uxn_c_l302_c2_9cba_return_output : unsigned(0 downto 0);

-- BIN_OP_GT[uxn_c_l311_c44_88dc]
signal BIN_OP_GT_uxn_c_l311_c44_88dc_left : unsigned(15 downto 0);
signal BIN_OP_GT_uxn_c_l311_c44_88dc_right : unsigned(15 downto 0);
signal BIN_OP_GT_uxn_c_l311_c44_88dc_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_c_l311_c65_3b56]
signal BIN_OP_PLUS_uxn_c_l311_c65_3b56_left : unsigned(23 downto 0);
signal BIN_OP_PLUS_uxn_c_l311_c65_3b56_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_c_l311_c65_3b56_return_output : unsigned(24 downto 0);

-- MUX[uxn_c_l311_c44_b965]
signal MUX_uxn_c_l311_c44_b965_cond : unsigned(0 downto 0);
signal MUX_uxn_c_l311_c44_b965_iftrue : unsigned(23 downto 0);
signal MUX_uxn_c_l311_c44_b965_iffalse : unsigned(23 downto 0);
signal MUX_uxn_c_l311_c44_b965_return_output : unsigned(23 downto 0);

-- MUX[uxn_c_l311_c16_5d3e]
signal MUX_uxn_c_l311_c16_5d3e_cond : unsigned(0 downto 0);
signal MUX_uxn_c_l311_c16_5d3e_iftrue : unsigned(23 downto 0);
signal MUX_uxn_c_l311_c16_5d3e_iffalse : unsigned(23 downto 0);
signal MUX_uxn_c_l311_c16_5d3e_return_output : unsigned(23 downto 0);

-- BIN_OP_EQ[uxn_c_l312_c16_4c21]
signal BIN_OP_EQ_uxn_c_l312_c16_4c21_left : unsigned(23 downto 0);
signal BIN_OP_EQ_uxn_c_l312_c16_4c21_right : unsigned(23 downto 0);
signal BIN_OP_EQ_uxn_c_l312_c16_4c21_return_output : unsigned(0 downto 0);

-- MUX[uxn_c_l312_c16_1944]
signal MUX_uxn_c_l312_c16_1944_cond : unsigned(0 downto 0);
signal MUX_uxn_c_l312_c16_1944_iftrue : unsigned(0 downto 0);
signal MUX_uxn_c_l312_c16_1944_iffalse : unsigned(0 downto 0);
signal MUX_uxn_c_l312_c16_1944_return_output : unsigned(0 downto 0);

-- MUX[uxn_c_l314_c16_61c4]
signal MUX_uxn_c_l314_c16_61c4_cond : unsigned(0 downto 0);
signal MUX_uxn_c_l314_c16_61c4_iftrue : unsigned(0 downto 0);
signal MUX_uxn_c_l314_c16_61c4_iffalse : unsigned(0 downto 0);
signal MUX_uxn_c_l314_c16_61c4_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_c_l314_c3_4639]
signal BIN_OP_PLUS_uxn_c_l314_c3_4639_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_c_l314_c3_4639_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_c_l314_c3_4639_return_output : unsigned(16 downto 0);

-- MUX[uxn_c_l315_c21_ddb1]
signal MUX_uxn_c_l315_c21_ddb1_cond : unsigned(0 downto 0);
signal MUX_uxn_c_l315_c21_ddb1_iftrue : unsigned(7 downto 0);
signal MUX_uxn_c_l315_c21_ddb1_iffalse : unsigned(7 downto 0);
signal MUX_uxn_c_l315_c21_ddb1_return_output : unsigned(7 downto 0);

-- UNARY_OP_NOT[uxn_c_l317_c14_2cfb]
signal UNARY_OP_NOT_uxn_c_l317_c14_2cfb_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_uxn_c_l317_c14_2cfb_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_c_l317_c1_20da]
signal TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_return_output : unsigned(0 downto 0);

-- u16_addr_MUX[uxn_c_l317_c9_9a0e]
signal u16_addr_MUX_uxn_c_l317_c9_9a0e_cond : unsigned(0 downto 0);
signal u16_addr_MUX_uxn_c_l317_c9_9a0e_iftrue : unsigned(15 downto 0);
signal u16_addr_MUX_uxn_c_l317_c9_9a0e_iffalse : unsigned(15 downto 0);
signal u16_addr_MUX_uxn_c_l317_c9_9a0e_return_output : unsigned(15 downto 0);

-- vram_write_layer_MUX[uxn_c_l317_c9_9a0e]
signal vram_write_layer_MUX_uxn_c_l317_c9_9a0e_cond : unsigned(0 downto 0);
signal vram_write_layer_MUX_uxn_c_l317_c9_9a0e_iftrue : unsigned(0 downto 0);
signal vram_write_layer_MUX_uxn_c_l317_c9_9a0e_iffalse : unsigned(0 downto 0);
signal vram_write_layer_MUX_uxn_c_l317_c9_9a0e_return_output : unsigned(0 downto 0);

-- device_ram_address_MUX[uxn_c_l317_c9_9a0e]
signal device_ram_address_MUX_uxn_c_l317_c9_9a0e_cond : unsigned(0 downto 0);
signal device_ram_address_MUX_uxn_c_l317_c9_9a0e_iftrue : unsigned(7 downto 0);
signal device_ram_address_MUX_uxn_c_l317_c9_9a0e_iffalse : unsigned(7 downto 0);
signal device_ram_address_MUX_uxn_c_l317_c9_9a0e_return_output : unsigned(7 downto 0);

-- is_device_ram_write_MUX[uxn_c_l317_c9_9a0e]
signal is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_cond : unsigned(0 downto 0);
signal is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_iftrue : unsigned(0 downto 0);
signal is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_iffalse : unsigned(0 downto 0);
signal is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_return_output : unsigned(0 downto 0);

-- is_ram_write_MUX[uxn_c_l317_c9_9a0e]
signal is_ram_write_MUX_uxn_c_l317_c9_9a0e_cond : unsigned(0 downto 0);
signal is_ram_write_MUX_uxn_c_l317_c9_9a0e_iftrue : unsigned(0 downto 0);
signal is_ram_write_MUX_uxn_c_l317_c9_9a0e_iffalse : unsigned(0 downto 0);
signal is_ram_write_MUX_uxn_c_l317_c9_9a0e_return_output : unsigned(0 downto 0);

-- is_vram_write_MUX[uxn_c_l317_c9_9a0e]
signal is_vram_write_MUX_uxn_c_l317_c9_9a0e_cond : unsigned(0 downto 0);
signal is_vram_write_MUX_uxn_c_l317_c9_9a0e_iftrue : unsigned(0 downto 0);
signal is_vram_write_MUX_uxn_c_l317_c9_9a0e_iffalse : unsigned(0 downto 0);
signal is_vram_write_MUX_uxn_c_l317_c9_9a0e_return_output : unsigned(0 downto 0);

-- vram_value_MUX[uxn_c_l317_c9_9a0e]
signal vram_value_MUX_uxn_c_l317_c9_9a0e_cond : unsigned(0 downto 0);
signal vram_value_MUX_uxn_c_l317_c9_9a0e_iftrue : unsigned(7 downto 0);
signal vram_value_MUX_uxn_c_l317_c9_9a0e_iffalse : unsigned(7 downto 0);
signal vram_value_MUX_uxn_c_l317_c9_9a0e_return_output : unsigned(7 downto 0);

-- ram_write_value_MUX[uxn_c_l317_c9_9a0e]
signal ram_write_value_MUX_uxn_c_l317_c9_9a0e_cond : unsigned(0 downto 0);
signal ram_write_value_MUX_uxn_c_l317_c9_9a0e_iftrue : unsigned(7 downto 0);
signal ram_write_value_MUX_uxn_c_l317_c9_9a0e_iffalse : unsigned(7 downto 0);
signal ram_write_value_MUX_uxn_c_l317_c9_9a0e_return_output : unsigned(7 downto 0);

-- cpu_step_result_MUX[uxn_c_l317_c9_9a0e]
signal cpu_step_result_MUX_uxn_c_l317_c9_9a0e_cond : unsigned(0 downto 0);
signal cpu_step_result_MUX_uxn_c_l317_c9_9a0e_iftrue : cpu_step_result_t;
signal cpu_step_result_MUX_uxn_c_l317_c9_9a0e_iffalse : cpu_step_result_t;
signal cpu_step_result_MUX_uxn_c_l317_c9_9a0e_return_output : cpu_step_result_t;

-- step_cpu[uxn_c_l318_c21_a9b6]
signal step_cpu_uxn_c_l318_c21_a9b6_CLOCK_ENABLE : unsigned(0 downto 0);
signal step_cpu_uxn_c_l318_c21_a9b6_previous_ram_read_value : unsigned(7 downto 0);
signal step_cpu_uxn_c_l318_c21_a9b6_previous_device_ram_read : unsigned(7 downto 0);
signal step_cpu_uxn_c_l318_c21_a9b6_use_vector : unsigned(0 downto 0);
signal step_cpu_uxn_c_l318_c21_a9b6_vector : unsigned(15 downto 0);
signal step_cpu_uxn_c_l318_c21_a9b6_return_output : cpu_step_result_t;

-- main_ram_update[uxn_c_l329_c19_6697]
signal main_ram_update_uxn_c_l329_c19_6697_CLOCK_ENABLE : unsigned(0 downto 0);
signal main_ram_update_uxn_c_l329_c19_6697_ram_address : unsigned(15 downto 0);
signal main_ram_update_uxn_c_l329_c19_6697_value : unsigned(7 downto 0);
signal main_ram_update_uxn_c_l329_c19_6697_write_enable : unsigned(0 downto 0);
signal main_ram_update_uxn_c_l329_c19_6697_return_output : unsigned(7 downto 0);

-- device_ram_update[uxn_c_l335_c26_db12]
signal device_ram_update_uxn_c_l335_c26_db12_CLOCK_ENABLE : unsigned(0 downto 0);
signal device_ram_update_uxn_c_l335_c26_db12_device_address : unsigned(7 downto 0);
signal device_ram_update_uxn_c_l335_c26_db12_value : unsigned(7 downto 0);
signal device_ram_update_uxn_c_l335_c26_db12_write_enable : unsigned(0 downto 0);
signal device_ram_update_uxn_c_l335_c26_db12_return_output : unsigned(7 downto 0);

-- step_gpu[uxn_c_l341_c20_9854]
signal step_gpu_uxn_c_l341_c20_9854_CLOCK_ENABLE : unsigned(0 downto 0);
signal step_gpu_uxn_c_l341_c20_9854_is_active_drawing_area : unsigned(0 downto 0);
signal step_gpu_uxn_c_l341_c20_9854_is_vram_write : unsigned(0 downto 0);
signal step_gpu_uxn_c_l341_c20_9854_vram_write_layer : unsigned(0 downto 0);
signal step_gpu_uxn_c_l341_c20_9854_vram_address : unsigned(15 downto 0);
signal step_gpu_uxn_c_l341_c20_9854_vram_value : unsigned(7 downto 0);
signal step_gpu_uxn_c_l341_c20_9854_return_output : gpu_step_result_t;

-- palette_snoop[uxn_c_l343_c20_f328]
signal palette_snoop_uxn_c_l343_c20_f328_CLOCK_ENABLE : unsigned(0 downto 0);
signal palette_snoop_uxn_c_l343_c20_f328_device_ram_address : unsigned(7 downto 0);
signal palette_snoop_uxn_c_l343_c20_f328_device_ram_value : unsigned(7 downto 0);
signal palette_snoop_uxn_c_l343_c20_f328_is_device_ram_write : unsigned(0 downto 0);
signal palette_snoop_uxn_c_l343_c20_f328_gpu_step_color : unsigned(1 downto 0);
signal palette_snoop_uxn_c_l343_c20_f328_return_output : unsigned(15 downto 0);

-- vector_snoop[uxn_c_l344_c18_80ab]
signal vector_snoop_uxn_c_l344_c18_80ab_CLOCK_ENABLE : unsigned(0 downto 0);
signal vector_snoop_uxn_c_l344_c18_80ab_device_ram_address : unsigned(7 downto 0);
signal vector_snoop_uxn_c_l344_c18_80ab_device_ram_value : unsigned(7 downto 0);
signal vector_snoop_uxn_c_l344_c18_80ab_is_device_ram_write : unsigned(0 downto 0);
signal vector_snoop_uxn_c_l344_c18_80ab_return_output : unsigned(15 downto 0);

-- BIN_OP_OR_uint1_t_uint1_t_uxn_c_l313_l314_DUPLICATE_e2dd
signal BIN_OP_OR_uint1_t_uint1_t_uxn_c_l313_l314_DUPLICATE_e2dd_left : unsigned(0 downto 0);
signal BIN_OP_OR_uint1_t_uint1_t_uxn_c_l313_l314_DUPLICATE_e2dd_right : unsigned(0 downto 0);
signal BIN_OP_OR_uint1_t_uint1_t_uxn_c_l313_l314_DUPLICATE_e2dd_return_output : unsigned(0 downto 0);


begin

-- SUBMODULE INSTANCES 
-- UNARY_OP_NOT_uxn_c_l302_c7_51e8
UNARY_OP_NOT_uxn_c_l302_c7_51e8 : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_uxn_c_l302_c7_51e8_expr,
UNARY_OP_NOT_uxn_c_l302_c7_51e8_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e
FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_return_output);

-- u16_addr_MUX_uxn_c_l302_c2_9cba
u16_addr_MUX_uxn_c_l302_c2_9cba : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
u16_addr_MUX_uxn_c_l302_c2_9cba_cond,
u16_addr_MUX_uxn_c_l302_c2_9cba_iftrue,
u16_addr_MUX_uxn_c_l302_c2_9cba_iffalse,
u16_addr_MUX_uxn_c_l302_c2_9cba_return_output);

-- vram_write_layer_MUX_uxn_c_l302_c2_9cba
vram_write_layer_MUX_uxn_c_l302_c2_9cba : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
vram_write_layer_MUX_uxn_c_l302_c2_9cba_cond,
vram_write_layer_MUX_uxn_c_l302_c2_9cba_iftrue,
vram_write_layer_MUX_uxn_c_l302_c2_9cba_iffalse,
vram_write_layer_MUX_uxn_c_l302_c2_9cba_return_output);

-- device_ram_address_MUX_uxn_c_l302_c2_9cba
device_ram_address_MUX_uxn_c_l302_c2_9cba : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
device_ram_address_MUX_uxn_c_l302_c2_9cba_cond,
device_ram_address_MUX_uxn_c_l302_c2_9cba_iftrue,
device_ram_address_MUX_uxn_c_l302_c2_9cba_iffalse,
device_ram_address_MUX_uxn_c_l302_c2_9cba_return_output);

-- is_device_ram_write_MUX_uxn_c_l302_c2_9cba
is_device_ram_write_MUX_uxn_c_l302_c2_9cba : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_device_ram_write_MUX_uxn_c_l302_c2_9cba_cond,
is_device_ram_write_MUX_uxn_c_l302_c2_9cba_iftrue,
is_device_ram_write_MUX_uxn_c_l302_c2_9cba_iffalse,
is_device_ram_write_MUX_uxn_c_l302_c2_9cba_return_output);

-- is_ram_write_MUX_uxn_c_l302_c2_9cba
is_ram_write_MUX_uxn_c_l302_c2_9cba : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_ram_write_MUX_uxn_c_l302_c2_9cba_cond,
is_ram_write_MUX_uxn_c_l302_c2_9cba_iftrue,
is_ram_write_MUX_uxn_c_l302_c2_9cba_iffalse,
is_ram_write_MUX_uxn_c_l302_c2_9cba_return_output);

-- is_vram_write_MUX_uxn_c_l302_c2_9cba
is_vram_write_MUX_uxn_c_l302_c2_9cba : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_vram_write_MUX_uxn_c_l302_c2_9cba_cond,
is_vram_write_MUX_uxn_c_l302_c2_9cba_iftrue,
is_vram_write_MUX_uxn_c_l302_c2_9cba_iffalse,
is_vram_write_MUX_uxn_c_l302_c2_9cba_return_output);

-- boot_check_MUX_uxn_c_l302_c2_9cba
boot_check_MUX_uxn_c_l302_c2_9cba : entity work.MUX_uint1_t_uint24_t_uint24_t_0CLK_de264c78 port map (
boot_check_MUX_uxn_c_l302_c2_9cba_cond,
boot_check_MUX_uxn_c_l302_c2_9cba_iftrue,
boot_check_MUX_uxn_c_l302_c2_9cba_iffalse,
boot_check_MUX_uxn_c_l302_c2_9cba_return_output);

-- vram_value_MUX_uxn_c_l302_c2_9cba
vram_value_MUX_uxn_c_l302_c2_9cba : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
vram_value_MUX_uxn_c_l302_c2_9cba_cond,
vram_value_MUX_uxn_c_l302_c2_9cba_iftrue,
vram_value_MUX_uxn_c_l302_c2_9cba_iffalse,
vram_value_MUX_uxn_c_l302_c2_9cba_return_output);

-- ram_write_value_MUX_uxn_c_l302_c2_9cba
ram_write_value_MUX_uxn_c_l302_c2_9cba : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ram_write_value_MUX_uxn_c_l302_c2_9cba_cond,
ram_write_value_MUX_uxn_c_l302_c2_9cba_iftrue,
ram_write_value_MUX_uxn_c_l302_c2_9cba_iffalse,
ram_write_value_MUX_uxn_c_l302_c2_9cba_return_output);

-- cpu_step_result_MUX_uxn_c_l302_c2_9cba
cpu_step_result_MUX_uxn_c_l302_c2_9cba : entity work.MUX_uint1_t_cpu_step_result_t_cpu_step_result_t_0CLK_de264c78 port map (
cpu_step_result_MUX_uxn_c_l302_c2_9cba_cond,
cpu_step_result_MUX_uxn_c_l302_c2_9cba_iftrue,
cpu_step_result_MUX_uxn_c_l302_c2_9cba_iffalse,
cpu_step_result_MUX_uxn_c_l302_c2_9cba_return_output);

-- is_booted_MUX_uxn_c_l302_c2_9cba
is_booted_MUX_uxn_c_l302_c2_9cba : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_booted_MUX_uxn_c_l302_c2_9cba_cond,
is_booted_MUX_uxn_c_l302_c2_9cba_iftrue,
is_booted_MUX_uxn_c_l302_c2_9cba_iffalse,
is_booted_MUX_uxn_c_l302_c2_9cba_return_output);

-- BIN_OP_GT_uxn_c_l311_c44_88dc
BIN_OP_GT_uxn_c_l311_c44_88dc : entity work.BIN_OP_GT_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_c_l311_c44_88dc_left,
BIN_OP_GT_uxn_c_l311_c44_88dc_right,
BIN_OP_GT_uxn_c_l311_c44_88dc_return_output);

-- BIN_OP_PLUS_uxn_c_l311_c65_3b56
BIN_OP_PLUS_uxn_c_l311_c65_3b56 : entity work.BIN_OP_PLUS_uint24_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_c_l311_c65_3b56_left,
BIN_OP_PLUS_uxn_c_l311_c65_3b56_right,
BIN_OP_PLUS_uxn_c_l311_c65_3b56_return_output);

-- MUX_uxn_c_l311_c44_b965
MUX_uxn_c_l311_c44_b965 : entity work.MUX_uint1_t_uint24_t_uint24_t_0CLK_de264c78 port map (
MUX_uxn_c_l311_c44_b965_cond,
MUX_uxn_c_l311_c44_b965_iftrue,
MUX_uxn_c_l311_c44_b965_iffalse,
MUX_uxn_c_l311_c44_b965_return_output);

-- MUX_uxn_c_l311_c16_5d3e
MUX_uxn_c_l311_c16_5d3e : entity work.MUX_uint1_t_uint24_t_uint24_t_0CLK_de264c78 port map (
MUX_uxn_c_l311_c16_5d3e_cond,
MUX_uxn_c_l311_c16_5d3e_iftrue,
MUX_uxn_c_l311_c16_5d3e_iffalse,
MUX_uxn_c_l311_c16_5d3e_return_output);

-- BIN_OP_EQ_uxn_c_l312_c16_4c21
BIN_OP_EQ_uxn_c_l312_c16_4c21 : entity work.BIN_OP_EQ_uint24_t_uint24_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_c_l312_c16_4c21_left,
BIN_OP_EQ_uxn_c_l312_c16_4c21_right,
BIN_OP_EQ_uxn_c_l312_c16_4c21_return_output);

-- MUX_uxn_c_l312_c16_1944
MUX_uxn_c_l312_c16_1944 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
MUX_uxn_c_l312_c16_1944_cond,
MUX_uxn_c_l312_c16_1944_iftrue,
MUX_uxn_c_l312_c16_1944_iffalse,
MUX_uxn_c_l312_c16_1944_return_output);

-- MUX_uxn_c_l314_c16_61c4
MUX_uxn_c_l314_c16_61c4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
MUX_uxn_c_l314_c16_61c4_cond,
MUX_uxn_c_l314_c16_61c4_iftrue,
MUX_uxn_c_l314_c16_61c4_iffalse,
MUX_uxn_c_l314_c16_61c4_return_output);

-- BIN_OP_PLUS_uxn_c_l314_c3_4639
BIN_OP_PLUS_uxn_c_l314_c3_4639 : entity work.BIN_OP_PLUS_uint16_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_c_l314_c3_4639_left,
BIN_OP_PLUS_uxn_c_l314_c3_4639_right,
BIN_OP_PLUS_uxn_c_l314_c3_4639_return_output);

-- MUX_uxn_c_l315_c21_ddb1
MUX_uxn_c_l315_c21_ddb1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_c_l315_c21_ddb1_cond,
MUX_uxn_c_l315_c21_ddb1_iftrue,
MUX_uxn_c_l315_c21_ddb1_iffalse,
MUX_uxn_c_l315_c21_ddb1_return_output);

-- UNARY_OP_NOT_uxn_c_l317_c14_2cfb
UNARY_OP_NOT_uxn_c_l317_c14_2cfb : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_uxn_c_l317_c14_2cfb_expr,
UNARY_OP_NOT_uxn_c_l317_c14_2cfb_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da
TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_return_output);

-- u16_addr_MUX_uxn_c_l317_c9_9a0e
u16_addr_MUX_uxn_c_l317_c9_9a0e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
u16_addr_MUX_uxn_c_l317_c9_9a0e_cond,
u16_addr_MUX_uxn_c_l317_c9_9a0e_iftrue,
u16_addr_MUX_uxn_c_l317_c9_9a0e_iffalse,
u16_addr_MUX_uxn_c_l317_c9_9a0e_return_output);

-- vram_write_layer_MUX_uxn_c_l317_c9_9a0e
vram_write_layer_MUX_uxn_c_l317_c9_9a0e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
vram_write_layer_MUX_uxn_c_l317_c9_9a0e_cond,
vram_write_layer_MUX_uxn_c_l317_c9_9a0e_iftrue,
vram_write_layer_MUX_uxn_c_l317_c9_9a0e_iffalse,
vram_write_layer_MUX_uxn_c_l317_c9_9a0e_return_output);

-- device_ram_address_MUX_uxn_c_l317_c9_9a0e
device_ram_address_MUX_uxn_c_l317_c9_9a0e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
device_ram_address_MUX_uxn_c_l317_c9_9a0e_cond,
device_ram_address_MUX_uxn_c_l317_c9_9a0e_iftrue,
device_ram_address_MUX_uxn_c_l317_c9_9a0e_iffalse,
device_ram_address_MUX_uxn_c_l317_c9_9a0e_return_output);

-- is_device_ram_write_MUX_uxn_c_l317_c9_9a0e
is_device_ram_write_MUX_uxn_c_l317_c9_9a0e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_cond,
is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_iftrue,
is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_iffalse,
is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_return_output);

-- is_ram_write_MUX_uxn_c_l317_c9_9a0e
is_ram_write_MUX_uxn_c_l317_c9_9a0e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_ram_write_MUX_uxn_c_l317_c9_9a0e_cond,
is_ram_write_MUX_uxn_c_l317_c9_9a0e_iftrue,
is_ram_write_MUX_uxn_c_l317_c9_9a0e_iffalse,
is_ram_write_MUX_uxn_c_l317_c9_9a0e_return_output);

-- is_vram_write_MUX_uxn_c_l317_c9_9a0e
is_vram_write_MUX_uxn_c_l317_c9_9a0e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_vram_write_MUX_uxn_c_l317_c9_9a0e_cond,
is_vram_write_MUX_uxn_c_l317_c9_9a0e_iftrue,
is_vram_write_MUX_uxn_c_l317_c9_9a0e_iffalse,
is_vram_write_MUX_uxn_c_l317_c9_9a0e_return_output);

-- vram_value_MUX_uxn_c_l317_c9_9a0e
vram_value_MUX_uxn_c_l317_c9_9a0e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
vram_value_MUX_uxn_c_l317_c9_9a0e_cond,
vram_value_MUX_uxn_c_l317_c9_9a0e_iftrue,
vram_value_MUX_uxn_c_l317_c9_9a0e_iffalse,
vram_value_MUX_uxn_c_l317_c9_9a0e_return_output);

-- ram_write_value_MUX_uxn_c_l317_c9_9a0e
ram_write_value_MUX_uxn_c_l317_c9_9a0e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ram_write_value_MUX_uxn_c_l317_c9_9a0e_cond,
ram_write_value_MUX_uxn_c_l317_c9_9a0e_iftrue,
ram_write_value_MUX_uxn_c_l317_c9_9a0e_iffalse,
ram_write_value_MUX_uxn_c_l317_c9_9a0e_return_output);

-- cpu_step_result_MUX_uxn_c_l317_c9_9a0e
cpu_step_result_MUX_uxn_c_l317_c9_9a0e : entity work.MUX_uint1_t_cpu_step_result_t_cpu_step_result_t_0CLK_de264c78 port map (
cpu_step_result_MUX_uxn_c_l317_c9_9a0e_cond,
cpu_step_result_MUX_uxn_c_l317_c9_9a0e_iftrue,
cpu_step_result_MUX_uxn_c_l317_c9_9a0e_iffalse,
cpu_step_result_MUX_uxn_c_l317_c9_9a0e_return_output);

-- step_cpu_uxn_c_l318_c21_a9b6
step_cpu_uxn_c_l318_c21_a9b6 : entity work.step_cpu_0CLK_d875878c port map (
clk,
step_cpu_uxn_c_l318_c21_a9b6_CLOCK_ENABLE,
step_cpu_uxn_c_l318_c21_a9b6_previous_ram_read_value,
step_cpu_uxn_c_l318_c21_a9b6_previous_device_ram_read,
step_cpu_uxn_c_l318_c21_a9b6_use_vector,
step_cpu_uxn_c_l318_c21_a9b6_vector,
step_cpu_uxn_c_l318_c21_a9b6_return_output);

-- main_ram_update_uxn_c_l329_c19_6697
main_ram_update_uxn_c_l329_c19_6697 : entity work.main_ram_update_0CLK_23f04728 port map (
clk,
main_ram_update_uxn_c_l329_c19_6697_CLOCK_ENABLE,
main_ram_update_uxn_c_l329_c19_6697_ram_address,
main_ram_update_uxn_c_l329_c19_6697_value,
main_ram_update_uxn_c_l329_c19_6697_write_enable,
main_ram_update_uxn_c_l329_c19_6697_return_output);

-- device_ram_update_uxn_c_l335_c26_db12
device_ram_update_uxn_c_l335_c26_db12 : entity work.device_ram_update_0CLK_23f04728 port map (
clk,
device_ram_update_uxn_c_l335_c26_db12_CLOCK_ENABLE,
device_ram_update_uxn_c_l335_c26_db12_device_address,
device_ram_update_uxn_c_l335_c26_db12_value,
device_ram_update_uxn_c_l335_c26_db12_write_enable,
device_ram_update_uxn_c_l335_c26_db12_return_output);

-- step_gpu_uxn_c_l341_c20_9854
step_gpu_uxn_c_l341_c20_9854 : entity work.step_gpu_0CLK_6d83165a port map (
clk,
step_gpu_uxn_c_l341_c20_9854_CLOCK_ENABLE,
step_gpu_uxn_c_l341_c20_9854_is_active_drawing_area,
step_gpu_uxn_c_l341_c20_9854_is_vram_write,
step_gpu_uxn_c_l341_c20_9854_vram_write_layer,
step_gpu_uxn_c_l341_c20_9854_vram_address,
step_gpu_uxn_c_l341_c20_9854_vram_value,
step_gpu_uxn_c_l341_c20_9854_return_output);

-- palette_snoop_uxn_c_l343_c20_f328
palette_snoop_uxn_c_l343_c20_f328 : entity work.palette_snoop_0CLK_ddbb7dc6 port map (
clk,
palette_snoop_uxn_c_l343_c20_f328_CLOCK_ENABLE,
palette_snoop_uxn_c_l343_c20_f328_device_ram_address,
palette_snoop_uxn_c_l343_c20_f328_device_ram_value,
palette_snoop_uxn_c_l343_c20_f328_is_device_ram_write,
palette_snoop_uxn_c_l343_c20_f328_gpu_step_color,
palette_snoop_uxn_c_l343_c20_f328_return_output);

-- vector_snoop_uxn_c_l344_c18_80ab
vector_snoop_uxn_c_l344_c18_80ab : entity work.vector_snoop_0CLK_10d8c973 port map (
clk,
vector_snoop_uxn_c_l344_c18_80ab_CLOCK_ENABLE,
vector_snoop_uxn_c_l344_c18_80ab_device_ram_address,
vector_snoop_uxn_c_l344_c18_80ab_device_ram_value,
vector_snoop_uxn_c_l344_c18_80ab_is_device_ram_write,
vector_snoop_uxn_c_l344_c18_80ab_return_output);

-- BIN_OP_OR_uint1_t_uint1_t_uxn_c_l313_l314_DUPLICATE_e2dd
BIN_OP_OR_uint1_t_uint1_t_uxn_c_l313_l314_DUPLICATE_e2dd : entity work.BIN_OP_OR_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_OR_uint1_t_uint1_t_uxn_c_l313_l314_DUPLICATE_e2dd_left,
BIN_OP_OR_uint1_t_uint1_t_uxn_c_l313_l314_DUPLICATE_e2dd_right,
BIN_OP_OR_uint1_t_uint1_t_uxn_c_l313_l314_DUPLICATE_e2dd_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 is_visible_pixel,
 rom_load_valid_byte,
 rom_load_address,
 rom_load_value,
 -- Registers
 boot_check,
 uxn_eval_result,
 is_booted,
 gpu_step_result,
 cpu_step_result,
 is_active_fill,
 is_ram_write,
 u16_addr,
 screen_vector,
 ram_write_value,
 ram_read_value,
 device_ram_address,
 device_ram_read_value,
 is_device_ram_write,
 is_vram_write,
 vram_write_layer,
 vram_value,
 -- All submodule outputs
 UNARY_OP_NOT_uxn_c_l302_c7_51e8_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_return_output,
 u16_addr_MUX_uxn_c_l302_c2_9cba_return_output,
 vram_write_layer_MUX_uxn_c_l302_c2_9cba_return_output,
 device_ram_address_MUX_uxn_c_l302_c2_9cba_return_output,
 is_device_ram_write_MUX_uxn_c_l302_c2_9cba_return_output,
 is_ram_write_MUX_uxn_c_l302_c2_9cba_return_output,
 is_vram_write_MUX_uxn_c_l302_c2_9cba_return_output,
 boot_check_MUX_uxn_c_l302_c2_9cba_return_output,
 vram_value_MUX_uxn_c_l302_c2_9cba_return_output,
 ram_write_value_MUX_uxn_c_l302_c2_9cba_return_output,
 cpu_step_result_MUX_uxn_c_l302_c2_9cba_return_output,
 is_booted_MUX_uxn_c_l302_c2_9cba_return_output,
 BIN_OP_GT_uxn_c_l311_c44_88dc_return_output,
 BIN_OP_PLUS_uxn_c_l311_c65_3b56_return_output,
 MUX_uxn_c_l311_c44_b965_return_output,
 MUX_uxn_c_l311_c16_5d3e_return_output,
 BIN_OP_EQ_uxn_c_l312_c16_4c21_return_output,
 MUX_uxn_c_l312_c16_1944_return_output,
 MUX_uxn_c_l314_c16_61c4_return_output,
 BIN_OP_PLUS_uxn_c_l314_c3_4639_return_output,
 MUX_uxn_c_l315_c21_ddb1_return_output,
 UNARY_OP_NOT_uxn_c_l317_c14_2cfb_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_return_output,
 u16_addr_MUX_uxn_c_l317_c9_9a0e_return_output,
 vram_write_layer_MUX_uxn_c_l317_c9_9a0e_return_output,
 device_ram_address_MUX_uxn_c_l317_c9_9a0e_return_output,
 is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_return_output,
 is_ram_write_MUX_uxn_c_l317_c9_9a0e_return_output,
 is_vram_write_MUX_uxn_c_l317_c9_9a0e_return_output,
 vram_value_MUX_uxn_c_l317_c9_9a0e_return_output,
 ram_write_value_MUX_uxn_c_l317_c9_9a0e_return_output,
 cpu_step_result_MUX_uxn_c_l317_c9_9a0e_return_output,
 step_cpu_uxn_c_l318_c21_a9b6_return_output,
 main_ram_update_uxn_c_l329_c19_6697_return_output,
 device_ram_update_uxn_c_l335_c26_db12_return_output,
 step_gpu_uxn_c_l341_c20_9854_return_output,
 palette_snoop_uxn_c_l343_c20_f328_return_output,
 vector_snoop_uxn_c_l344_c18_80ab_return_output,
 BIN_OP_OR_uint1_t_uint1_t_uxn_c_l313_l314_DUPLICATE_e2dd_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(15 downto 0);
 variable VAR_is_visible_pixel : unsigned(0 downto 0);
 variable VAR_rom_load_valid_byte : unsigned(0 downto 0);
 variable VAR_rom_load_address : unsigned(15 downto 0);
 variable VAR_rom_load_value : unsigned(7 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_c_l302_c7_51e8_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_c_l302_c7_51e8_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_iffalse : unsigned(0 downto 0);
 variable VAR_u16_addr_MUX_uxn_c_l302_c2_9cba_iftrue : unsigned(15 downto 0);
 variable VAR_u16_addr_uxn_c_l314_c3_4336 : unsigned(15 downto 0);
 variable VAR_u16_addr_MUX_uxn_c_l302_c2_9cba_iffalse : unsigned(15 downto 0);
 variable VAR_u16_addr_MUX_uxn_c_l317_c9_9a0e_return_output : unsigned(15 downto 0);
 variable VAR_u16_addr_MUX_uxn_c_l302_c2_9cba_return_output : unsigned(15 downto 0);
 variable VAR_u16_addr_MUX_uxn_c_l302_c2_9cba_cond : unsigned(0 downto 0);
 variable VAR_vram_write_layer_MUX_uxn_c_l302_c2_9cba_iftrue : unsigned(0 downto 0);
 variable VAR_vram_write_layer_MUX_uxn_c_l302_c2_9cba_iffalse : unsigned(0 downto 0);
 variable VAR_vram_write_layer_MUX_uxn_c_l317_c9_9a0e_return_output : unsigned(0 downto 0);
 variable VAR_vram_write_layer_MUX_uxn_c_l302_c2_9cba_return_output : unsigned(0 downto 0);
 variable VAR_vram_write_layer_MUX_uxn_c_l302_c2_9cba_cond : unsigned(0 downto 0);
 variable VAR_device_ram_address_MUX_uxn_c_l302_c2_9cba_iftrue : unsigned(7 downto 0);
 variable VAR_device_ram_address_MUX_uxn_c_l302_c2_9cba_iffalse : unsigned(7 downto 0);
 variable VAR_device_ram_address_MUX_uxn_c_l317_c9_9a0e_return_output : unsigned(7 downto 0);
 variable VAR_device_ram_address_MUX_uxn_c_l302_c2_9cba_return_output : unsigned(7 downto 0);
 variable VAR_device_ram_address_MUX_uxn_c_l302_c2_9cba_cond : unsigned(0 downto 0);
 variable VAR_is_device_ram_write_MUX_uxn_c_l302_c2_9cba_iftrue : unsigned(0 downto 0);
 variable VAR_is_device_ram_write_MUX_uxn_c_l302_c2_9cba_iffalse : unsigned(0 downto 0);
 variable VAR_is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_return_output : unsigned(0 downto 0);
 variable VAR_is_device_ram_write_MUX_uxn_c_l302_c2_9cba_return_output : unsigned(0 downto 0);
 variable VAR_is_device_ram_write_MUX_uxn_c_l302_c2_9cba_cond : unsigned(0 downto 0);
 variable VAR_is_ram_write_MUX_uxn_c_l302_c2_9cba_iftrue : unsigned(0 downto 0);
 variable VAR_is_ram_write_MUX_uxn_c_l302_c2_9cba_iffalse : unsigned(0 downto 0);
 variable VAR_is_ram_write_MUX_uxn_c_l317_c9_9a0e_return_output : unsigned(0 downto 0);
 variable VAR_is_ram_write_MUX_uxn_c_l302_c2_9cba_return_output : unsigned(0 downto 0);
 variable VAR_is_ram_write_MUX_uxn_c_l302_c2_9cba_cond : unsigned(0 downto 0);
 variable VAR_is_vram_write_MUX_uxn_c_l302_c2_9cba_iftrue : unsigned(0 downto 0);
 variable VAR_is_vram_write_MUX_uxn_c_l302_c2_9cba_iffalse : unsigned(0 downto 0);
 variable VAR_is_vram_write_MUX_uxn_c_l317_c9_9a0e_return_output : unsigned(0 downto 0);
 variable VAR_is_vram_write_MUX_uxn_c_l302_c2_9cba_return_output : unsigned(0 downto 0);
 variable VAR_is_vram_write_MUX_uxn_c_l302_c2_9cba_cond : unsigned(0 downto 0);
 variable VAR_boot_check_MUX_uxn_c_l302_c2_9cba_iftrue : unsigned(23 downto 0);
 variable VAR_boot_check_MUX_uxn_c_l302_c2_9cba_iffalse : unsigned(23 downto 0);
 variable VAR_boot_check_MUX_uxn_c_l302_c2_9cba_return_output : unsigned(23 downto 0);
 variable VAR_boot_check_MUX_uxn_c_l302_c2_9cba_cond : unsigned(0 downto 0);
 variable VAR_vram_value_MUX_uxn_c_l302_c2_9cba_iftrue : unsigned(7 downto 0);
 variable VAR_vram_value_MUX_uxn_c_l302_c2_9cba_iffalse : unsigned(7 downto 0);
 variable VAR_vram_value_MUX_uxn_c_l317_c9_9a0e_return_output : unsigned(7 downto 0);
 variable VAR_vram_value_MUX_uxn_c_l302_c2_9cba_return_output : unsigned(7 downto 0);
 variable VAR_vram_value_MUX_uxn_c_l302_c2_9cba_cond : unsigned(0 downto 0);
 variable VAR_ram_write_value_MUX_uxn_c_l302_c2_9cba_iftrue : unsigned(7 downto 0);
 variable VAR_ram_write_value_MUX_uxn_c_l302_c2_9cba_iffalse : unsigned(7 downto 0);
 variable VAR_ram_write_value_MUX_uxn_c_l317_c9_9a0e_return_output : unsigned(7 downto 0);
 variable VAR_ram_write_value_MUX_uxn_c_l302_c2_9cba_return_output : unsigned(7 downto 0);
 variable VAR_ram_write_value_MUX_uxn_c_l302_c2_9cba_cond : unsigned(0 downto 0);
 variable VAR_cpu_step_result_MUX_uxn_c_l302_c2_9cba_iftrue : cpu_step_result_t;
 variable VAR_cpu_step_result_MUX_uxn_c_l302_c2_9cba_iffalse : cpu_step_result_t;
 variable VAR_cpu_step_result_MUX_uxn_c_l317_c9_9a0e_return_output : cpu_step_result_t;
 variable VAR_cpu_step_result_MUX_uxn_c_l302_c2_9cba_return_output : cpu_step_result_t;
 variable VAR_cpu_step_result_MUX_uxn_c_l302_c2_9cba_cond : unsigned(0 downto 0);
 variable VAR_is_booted_MUX_uxn_c_l302_c2_9cba_iftrue : unsigned(0 downto 0);
 variable VAR_is_booted_MUX_uxn_c_l302_c2_9cba_iffalse : unsigned(0 downto 0);
 variable VAR_is_booted_MUX_uxn_c_l302_c2_9cba_return_output : unsigned(0 downto 0);
 variable VAR_is_booted_MUX_uxn_c_l302_c2_9cba_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_c_l311_c16_5d3e_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_c_l311_c16_5d3e_iftrue : unsigned(23 downto 0);
 variable VAR_MUX_uxn_c_l311_c16_5d3e_iffalse : unsigned(23 downto 0);
 variable VAR_MUX_uxn_c_l311_c44_b965_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_c_l311_c44_88dc_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_GT_uxn_c_l311_c44_88dc_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_GT_uxn_c_l311_c44_88dc_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_c_l311_c44_b965_iftrue : unsigned(23 downto 0);
 variable VAR_MUX_uxn_c_l311_c44_b965_iffalse : unsigned(23 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_c_l311_c65_3b56_left : unsigned(23 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_c_l311_c65_3b56_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_c_l311_c65_3b56_return_output : unsigned(24 downto 0);
 variable VAR_MUX_uxn_c_l311_c44_b965_return_output : unsigned(23 downto 0);
 variable VAR_MUX_uxn_c_l311_c16_5d3e_return_output : unsigned(23 downto 0);
 variable VAR_MUX_uxn_c_l312_c16_1944_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_c_l312_c16_4c21_left : unsigned(23 downto 0);
 variable VAR_BIN_OP_EQ_uxn_c_l312_c16_4c21_right : unsigned(23 downto 0);
 variable VAR_BIN_OP_EQ_uxn_c_l312_c16_4c21_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_c_l312_c16_1944_iftrue : unsigned(0 downto 0);
 variable VAR_MUX_uxn_c_l312_c16_1944_iffalse : unsigned(0 downto 0);
 variable VAR_MUX_uxn_c_l312_c16_1944_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_c_l314_c3_4639_left : unsigned(15 downto 0);
 variable VAR_MUX_uxn_c_l314_c16_61c4_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_c_l314_c16_61c4_iftrue : unsigned(0 downto 0);
 variable VAR_MUX_uxn_c_l314_c16_61c4_iffalse : unsigned(0 downto 0);
 variable VAR_MUX_uxn_c_l314_c16_61c4_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_c_l314_c3_4639_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_c_l314_c3_4639_return_output : unsigned(16 downto 0);
 variable VAR_MUX_uxn_c_l315_c21_ddb1_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_c_l315_c21_ddb1_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_c_l315_c21_ddb1_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_c_l315_c21_ddb1_return_output : unsigned(7 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_c_l317_c14_2cfb_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_c_l317_c14_2cfb_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_iffalse : unsigned(0 downto 0);
 variable VAR_u16_addr_MUX_uxn_c_l317_c9_9a0e_iftrue : unsigned(15 downto 0);
 variable VAR_u16_addr_MUX_uxn_c_l317_c9_9a0e_iffalse : unsigned(15 downto 0);
 variable VAR_u16_addr_MUX_uxn_c_l317_c9_9a0e_cond : unsigned(0 downto 0);
 variable VAR_vram_write_layer_MUX_uxn_c_l317_c9_9a0e_iftrue : unsigned(0 downto 0);
 variable VAR_vram_write_layer_MUX_uxn_c_l317_c9_9a0e_iffalse : unsigned(0 downto 0);
 variable VAR_vram_write_layer_MUX_uxn_c_l317_c9_9a0e_cond : unsigned(0 downto 0);
 variable VAR_device_ram_address_MUX_uxn_c_l317_c9_9a0e_iftrue : unsigned(7 downto 0);
 variable VAR_device_ram_address_MUX_uxn_c_l317_c9_9a0e_iffalse : unsigned(7 downto 0);
 variable VAR_device_ram_address_MUX_uxn_c_l317_c9_9a0e_cond : unsigned(0 downto 0);
 variable VAR_is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_iftrue : unsigned(0 downto 0);
 variable VAR_is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_iffalse : unsigned(0 downto 0);
 variable VAR_is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_cond : unsigned(0 downto 0);
 variable VAR_is_ram_write_MUX_uxn_c_l317_c9_9a0e_iftrue : unsigned(0 downto 0);
 variable VAR_is_ram_write_MUX_uxn_c_l317_c9_9a0e_iffalse : unsigned(0 downto 0);
 variable VAR_is_ram_write_MUX_uxn_c_l317_c9_9a0e_cond : unsigned(0 downto 0);
 variable VAR_is_vram_write_MUX_uxn_c_l317_c9_9a0e_iftrue : unsigned(0 downto 0);
 variable VAR_is_vram_write_MUX_uxn_c_l317_c9_9a0e_iffalse : unsigned(0 downto 0);
 variable VAR_is_vram_write_MUX_uxn_c_l317_c9_9a0e_cond : unsigned(0 downto 0);
 variable VAR_vram_value_MUX_uxn_c_l317_c9_9a0e_iftrue : unsigned(7 downto 0);
 variable VAR_vram_value_MUX_uxn_c_l317_c9_9a0e_iffalse : unsigned(7 downto 0);
 variable VAR_vram_value_MUX_uxn_c_l317_c9_9a0e_cond : unsigned(0 downto 0);
 variable VAR_ram_write_value_MUX_uxn_c_l317_c9_9a0e_iftrue : unsigned(7 downto 0);
 variable VAR_ram_write_value_MUX_uxn_c_l317_c9_9a0e_iffalse : unsigned(7 downto 0);
 variable VAR_ram_write_value_MUX_uxn_c_l317_c9_9a0e_cond : unsigned(0 downto 0);
 variable VAR_cpu_step_result_MUX_uxn_c_l317_c9_9a0e_iftrue : cpu_step_result_t;
 variable VAR_cpu_step_result_MUX_uxn_c_l317_c9_9a0e_iffalse : cpu_step_result_t;
 variable VAR_cpu_step_result_MUX_uxn_c_l317_c9_9a0e_cond : unsigned(0 downto 0);
 variable VAR_step_cpu_uxn_c_l318_c21_a9b6_previous_ram_read_value : unsigned(7 downto 0);
 variable VAR_step_cpu_uxn_c_l318_c21_a9b6_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_step_cpu_uxn_c_l318_c21_a9b6_use_vector : unsigned(0 downto 0);
 variable VAR_step_cpu_uxn_c_l318_c21_a9b6_vector : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_gpu_step_result_t_is_new_frame_d41d_uxn_c_l318_c69_6e2d_return_output : unsigned(0 downto 0);
 variable VAR_step_cpu_uxn_c_l318_c21_a9b6_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_step_cpu_uxn_c_l318_c21_a9b6_return_output : cpu_step_result_t;
 variable VAR_CONST_REF_RD_uint1_t_cpu_step_result_t_is_ram_write_d41d_uxn_c_l319_c18_e6d8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_cpu_step_result_t_u16_addr_d41d_uxn_c_l320_c14_8d49_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_cpu_step_result_t_device_ram_address_d41d_uxn_c_l321_c24_5ea8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_cpu_step_result_t_is_device_ram_write_d41d_uxn_c_l322_c25_df61_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_cpu_step_result_t_is_vram_write_d41d_uxn_c_l324_c19_bd0b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_cpu_step_result_t_vram_write_layer_d41d_uxn_c_l325_c22_9ead_return_output : unsigned(0 downto 0);
 variable VAR_main_ram_update_uxn_c_l329_c19_6697_ram_address : unsigned(15 downto 0);
 variable VAR_main_ram_update_uxn_c_l329_c19_6697_value : unsigned(7 downto 0);
 variable VAR_main_ram_update_uxn_c_l329_c19_6697_write_enable : unsigned(0 downto 0);
 variable VAR_main_ram_update_uxn_c_l329_c19_6697_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_main_ram_update_uxn_c_l329_c19_6697_return_output : unsigned(7 downto 0);
 variable VAR_device_ram_update_uxn_c_l335_c26_db12_device_address : unsigned(7 downto 0);
 variable VAR_device_ram_update_uxn_c_l335_c26_db12_value : unsigned(7 downto 0);
 variable VAR_device_ram_update_uxn_c_l335_c26_db12_write_enable : unsigned(0 downto 0);
 variable VAR_device_ram_update_uxn_c_l335_c26_db12_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_device_ram_update_uxn_c_l335_c26_db12_return_output : unsigned(7 downto 0);
 variable VAR_step_gpu_uxn_c_l341_c20_9854_is_active_drawing_area : unsigned(0 downto 0);
 variable VAR_step_gpu_uxn_c_l341_c20_9854_is_vram_write : unsigned(0 downto 0);
 variable VAR_step_gpu_uxn_c_l341_c20_9854_vram_write_layer : unsigned(0 downto 0);
 variable VAR_step_gpu_uxn_c_l341_c20_9854_vram_address : unsigned(15 downto 0);
 variable VAR_step_gpu_uxn_c_l341_c20_9854_vram_value : unsigned(7 downto 0);
 variable VAR_step_gpu_uxn_c_l341_c20_9854_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_step_gpu_uxn_c_l341_c20_9854_return_output : gpu_step_result_t;
 variable VAR_CONST_REF_RD_uint1_t_gpu_step_result_t_is_active_fill_d41d_uxn_c_l342_c19_b60d_return_output : unsigned(0 downto 0);
 variable VAR_palette_snoop_uxn_c_l343_c20_f328_device_ram_address : unsigned(7 downto 0);
 variable VAR_palette_snoop_uxn_c_l343_c20_f328_device_ram_value : unsigned(7 downto 0);
 variable VAR_palette_snoop_uxn_c_l343_c20_f328_is_device_ram_write : unsigned(0 downto 0);
 variable VAR_palette_snoop_uxn_c_l343_c20_f328_gpu_step_color : unsigned(1 downto 0);
 variable VAR_CONST_REF_RD_uint2_t_gpu_step_result_t_color_d41d_uxn_c_l343_c92_ec5c_return_output : unsigned(1 downto 0);
 variable VAR_palette_snoop_uxn_c_l343_c20_f328_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_palette_snoop_uxn_c_l343_c20_f328_return_output : unsigned(15 downto 0);
 variable VAR_vector_snoop_uxn_c_l344_c18_80ab_device_ram_address : unsigned(7 downto 0);
 variable VAR_vector_snoop_uxn_c_l344_c18_80ab_device_ram_value : unsigned(7 downto 0);
 variable VAR_vector_snoop_uxn_c_l344_c18_80ab_is_device_ram_write : unsigned(0 downto 0);
 variable VAR_vector_snoop_uxn_c_l344_c18_80ab_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_vector_snoop_uxn_c_l344_c18_80ab_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uint1_t_uint1_t_uxn_c_l313_l314_DUPLICATE_e2dd_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uint1_t_uint1_t_uxn_c_l313_l314_DUPLICATE_e2dd_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uint1_t_uint1_t_uxn_c_l313_l314_DUPLICATE_e2dd_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_cpu_step_result_t_u8_value_d41d_uxn_c_l323_l326_DUPLICATE_30f9_return_output : unsigned(7 downto 0);
 -- State registers comb logic variables
variable REG_VAR_boot_check : unsigned(23 downto 0);
variable REG_VAR_uxn_eval_result : unsigned(15 downto 0);
variable REG_VAR_is_booted : unsigned(0 downto 0);
variable REG_VAR_gpu_step_result : gpu_step_result_t;
variable REG_VAR_cpu_step_result : cpu_step_result_t;
variable REG_VAR_is_active_fill : unsigned(0 downto 0);
variable REG_VAR_is_ram_write : unsigned(0 downto 0);
variable REG_VAR_u16_addr : unsigned(15 downto 0);
variable REG_VAR_screen_vector : unsigned(15 downto 0);
variable REG_VAR_ram_write_value : unsigned(7 downto 0);
variable REG_VAR_ram_read_value : unsigned(7 downto 0);
variable REG_VAR_device_ram_address : unsigned(7 downto 0);
variable REG_VAR_device_ram_read_value : unsigned(7 downto 0);
variable REG_VAR_is_device_ram_write : unsigned(0 downto 0);
variable REG_VAR_is_vram_write : unsigned(0 downto 0);
variable REG_VAR_vram_write_layer : unsigned(0 downto 0);
variable REG_VAR_vram_value : unsigned(7 downto 0);
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_boot_check := boot_check;
  REG_VAR_uxn_eval_result := uxn_eval_result;
  REG_VAR_is_booted := is_booted;
  REG_VAR_gpu_step_result := gpu_step_result;
  REG_VAR_cpu_step_result := cpu_step_result;
  REG_VAR_is_active_fill := is_active_fill;
  REG_VAR_is_ram_write := is_ram_write;
  REG_VAR_u16_addr := u16_addr;
  REG_VAR_screen_vector := screen_vector;
  REG_VAR_ram_write_value := ram_write_value;
  REG_VAR_ram_read_value := ram_read_value;
  REG_VAR_device_ram_address := device_ram_address;
  REG_VAR_device_ram_read_value := device_ram_read_value;
  REG_VAR_is_device_ram_write := is_device_ram_write;
  REG_VAR_is_vram_write := is_vram_write;
  REG_VAR_vram_write_layer := vram_write_layer;
  REG_VAR_vram_value := vram_value;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_MUX_uxn_c_l314_c16_61c4_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_c_l312_c16_4c21_right := to_unsigned(16777215, 24);
     VAR_MUX_uxn_c_l314_c16_61c4_iffalse := to_unsigned(0, 1);
     VAR_MUX_uxn_c_l312_c16_1944_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_c_l312_c16_1944_iffalse := to_unsigned(0, 1);
     VAR_MUX_uxn_c_l311_c16_5d3e_iftrue := resize(to_unsigned(0, 1), 24);
     VAR_MUX_uxn_c_l311_c44_b965_iffalse := resize(to_unsigned(0, 1), 24);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_GT_uxn_c_l311_c44_88dc_right := to_unsigned(255, 16);
     VAR_BIN_OP_PLUS_uxn_c_l311_c65_3b56_right := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_iffalse := to_unsigned(0, 1);
     VAR_MUX_uxn_c_l315_c21_ddb1_iftrue := resize(to_unsigned(0, 1), 8);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_is_visible_pixel := is_visible_pixel;
     VAR_rom_load_valid_byte := rom_load_valid_byte;
     VAR_rom_load_address := rom_load_address;
     VAR_rom_load_value := rom_load_value;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_iffalse := VAR_CLOCK_ENABLE;
     VAR_device_ram_update_uxn_c_l335_c26_db12_CLOCK_ENABLE := VAR_CLOCK_ENABLE;
     VAR_main_ram_update_uxn_c_l329_c19_6697_CLOCK_ENABLE := VAR_CLOCK_ENABLE;
     VAR_palette_snoop_uxn_c_l343_c20_f328_CLOCK_ENABLE := VAR_CLOCK_ENABLE;
     VAR_step_gpu_uxn_c_l341_c20_9854_CLOCK_ENABLE := VAR_CLOCK_ENABLE;
     VAR_vector_snoop_uxn_c_l344_c18_80ab_CLOCK_ENABLE := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_PLUS_uxn_c_l311_c65_3b56_left := boot_check;
     VAR_boot_check_MUX_uxn_c_l302_c2_9cba_iffalse := boot_check;
     VAR_cpu_step_result_MUX_uxn_c_l302_c2_9cba_iftrue := cpu_step_result;
     VAR_cpu_step_result_MUX_uxn_c_l317_c9_9a0e_iffalse := cpu_step_result;
     VAR_device_ram_address_MUX_uxn_c_l302_c2_9cba_iftrue := device_ram_address;
     VAR_device_ram_address_MUX_uxn_c_l317_c9_9a0e_iffalse := device_ram_address;
     VAR_step_cpu_uxn_c_l318_c21_a9b6_previous_device_ram_read := device_ram_read_value;
     VAR_UNARY_OP_NOT_uxn_c_l317_c14_2cfb_expr := is_active_fill;
     VAR_UNARY_OP_NOT_uxn_c_l302_c7_51e8_expr := is_booted;
     VAR_is_booted_MUX_uxn_c_l302_c2_9cba_iffalse := is_booted;
     VAR_is_device_ram_write_MUX_uxn_c_l302_c2_9cba_iftrue := is_device_ram_write;
     VAR_is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_iffalse := is_device_ram_write;
     VAR_is_ram_write_MUX_uxn_c_l317_c9_9a0e_iffalse := is_ram_write;
     VAR_step_gpu_uxn_c_l341_c20_9854_is_active_drawing_area := VAR_is_visible_pixel;
     VAR_is_vram_write_MUX_uxn_c_l302_c2_9cba_iftrue := is_vram_write;
     VAR_is_vram_write_MUX_uxn_c_l317_c9_9a0e_iffalse := is_vram_write;
     VAR_step_cpu_uxn_c_l318_c21_a9b6_previous_ram_read_value := ram_read_value;
     VAR_ram_write_value_MUX_uxn_c_l317_c9_9a0e_iffalse := ram_write_value;
     VAR_BIN_OP_OR_uint1_t_uint1_t_uxn_c_l313_l314_DUPLICATE_e2dd_left := VAR_rom_load_valid_byte;
     VAR_MUX_uxn_c_l311_c16_5d3e_cond := VAR_rom_load_valid_byte;
     VAR_MUX_uxn_c_l315_c21_ddb1_iffalse := VAR_rom_load_value;
     VAR_step_cpu_uxn_c_l318_c21_a9b6_vector := screen_vector;
     VAR_BIN_OP_GT_uxn_c_l311_c44_88dc_left := u16_addr;
     VAR_BIN_OP_PLUS_uxn_c_l314_c3_4639_left := u16_addr;
     VAR_u16_addr_MUX_uxn_c_l317_c9_9a0e_iffalse := u16_addr;
     VAR_vram_value_MUX_uxn_c_l302_c2_9cba_iftrue := vram_value;
     VAR_vram_value_MUX_uxn_c_l317_c9_9a0e_iffalse := vram_value;
     VAR_vram_write_layer_MUX_uxn_c_l302_c2_9cba_iftrue := vram_write_layer;
     VAR_vram_write_layer_MUX_uxn_c_l317_c9_9a0e_iffalse := vram_write_layer;
     -- BIN_OP_GT[uxn_c_l311_c44_88dc] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_c_l311_c44_88dc_left <= VAR_BIN_OP_GT_uxn_c_l311_c44_88dc_left;
     BIN_OP_GT_uxn_c_l311_c44_88dc_right <= VAR_BIN_OP_GT_uxn_c_l311_c44_88dc_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_c_l311_c44_88dc_return_output := BIN_OP_GT_uxn_c_l311_c44_88dc_return_output;

     -- BIN_OP_PLUS[uxn_c_l311_c65_3b56] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_c_l311_c65_3b56_left <= VAR_BIN_OP_PLUS_uxn_c_l311_c65_3b56_left;
     BIN_OP_PLUS_uxn_c_l311_c65_3b56_right <= VAR_BIN_OP_PLUS_uxn_c_l311_c65_3b56_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_c_l311_c65_3b56_return_output := BIN_OP_PLUS_uxn_c_l311_c65_3b56_return_output;

     -- UNARY_OP_NOT[uxn_c_l317_c14_2cfb] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_uxn_c_l317_c14_2cfb_expr <= VAR_UNARY_OP_NOT_uxn_c_l317_c14_2cfb_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_uxn_c_l317_c14_2cfb_return_output := UNARY_OP_NOT_uxn_c_l317_c14_2cfb_return_output;

     -- CONST_REF_RD_uint1_t_gpu_step_result_t_is_new_frame_d41d[uxn_c_l318_c69_6e2d] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_gpu_step_result_t_is_new_frame_d41d_uxn_c_l318_c69_6e2d_return_output := gpu_step_result.is_new_frame;

     -- UNARY_OP_NOT[uxn_c_l302_c7_51e8] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_uxn_c_l302_c7_51e8_expr <= VAR_UNARY_OP_NOT_uxn_c_l302_c7_51e8_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_uxn_c_l302_c7_51e8_return_output := UNARY_OP_NOT_uxn_c_l302_c7_51e8_return_output;

     -- Submodule level 1
     VAR_MUX_uxn_c_l311_c44_b965_cond := VAR_BIN_OP_GT_uxn_c_l311_c44_88dc_return_output;
     VAR_MUX_uxn_c_l311_c44_b965_iftrue := resize(VAR_BIN_OP_PLUS_uxn_c_l311_c65_3b56_return_output, 24);
     VAR_step_cpu_uxn_c_l318_c21_a9b6_use_vector := VAR_CONST_REF_RD_uint1_t_gpu_step_result_t_is_new_frame_d41d_uxn_c_l318_c69_6e2d_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_cond := VAR_UNARY_OP_NOT_uxn_c_l302_c7_51e8_return_output;
     VAR_boot_check_MUX_uxn_c_l302_c2_9cba_cond := VAR_UNARY_OP_NOT_uxn_c_l302_c7_51e8_return_output;
     VAR_cpu_step_result_MUX_uxn_c_l302_c2_9cba_cond := VAR_UNARY_OP_NOT_uxn_c_l302_c7_51e8_return_output;
     VAR_device_ram_address_MUX_uxn_c_l302_c2_9cba_cond := VAR_UNARY_OP_NOT_uxn_c_l302_c7_51e8_return_output;
     VAR_is_booted_MUX_uxn_c_l302_c2_9cba_cond := VAR_UNARY_OP_NOT_uxn_c_l302_c7_51e8_return_output;
     VAR_is_device_ram_write_MUX_uxn_c_l302_c2_9cba_cond := VAR_UNARY_OP_NOT_uxn_c_l302_c7_51e8_return_output;
     VAR_is_ram_write_MUX_uxn_c_l302_c2_9cba_cond := VAR_UNARY_OP_NOT_uxn_c_l302_c7_51e8_return_output;
     VAR_is_vram_write_MUX_uxn_c_l302_c2_9cba_cond := VAR_UNARY_OP_NOT_uxn_c_l302_c7_51e8_return_output;
     VAR_ram_write_value_MUX_uxn_c_l302_c2_9cba_cond := VAR_UNARY_OP_NOT_uxn_c_l302_c7_51e8_return_output;
     VAR_u16_addr_MUX_uxn_c_l302_c2_9cba_cond := VAR_UNARY_OP_NOT_uxn_c_l302_c7_51e8_return_output;
     VAR_vram_value_MUX_uxn_c_l302_c2_9cba_cond := VAR_UNARY_OP_NOT_uxn_c_l302_c7_51e8_return_output;
     VAR_vram_write_layer_MUX_uxn_c_l302_c2_9cba_cond := VAR_UNARY_OP_NOT_uxn_c_l302_c7_51e8_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_cond := VAR_UNARY_OP_NOT_uxn_c_l317_c14_2cfb_return_output;
     VAR_cpu_step_result_MUX_uxn_c_l317_c9_9a0e_cond := VAR_UNARY_OP_NOT_uxn_c_l317_c14_2cfb_return_output;
     VAR_device_ram_address_MUX_uxn_c_l317_c9_9a0e_cond := VAR_UNARY_OP_NOT_uxn_c_l317_c14_2cfb_return_output;
     VAR_is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_cond := VAR_UNARY_OP_NOT_uxn_c_l317_c14_2cfb_return_output;
     VAR_is_ram_write_MUX_uxn_c_l317_c9_9a0e_cond := VAR_UNARY_OP_NOT_uxn_c_l317_c14_2cfb_return_output;
     VAR_is_vram_write_MUX_uxn_c_l317_c9_9a0e_cond := VAR_UNARY_OP_NOT_uxn_c_l317_c14_2cfb_return_output;
     VAR_ram_write_value_MUX_uxn_c_l317_c9_9a0e_cond := VAR_UNARY_OP_NOT_uxn_c_l317_c14_2cfb_return_output;
     VAR_u16_addr_MUX_uxn_c_l317_c9_9a0e_cond := VAR_UNARY_OP_NOT_uxn_c_l317_c14_2cfb_return_output;
     VAR_vram_value_MUX_uxn_c_l317_c9_9a0e_cond := VAR_UNARY_OP_NOT_uxn_c_l317_c14_2cfb_return_output;
     VAR_vram_write_layer_MUX_uxn_c_l317_c9_9a0e_cond := VAR_UNARY_OP_NOT_uxn_c_l317_c14_2cfb_return_output;
     -- MUX[uxn_c_l311_c44_b965] LATENCY=0
     -- Inputs
     MUX_uxn_c_l311_c44_b965_cond <= VAR_MUX_uxn_c_l311_c44_b965_cond;
     MUX_uxn_c_l311_c44_b965_iftrue <= VAR_MUX_uxn_c_l311_c44_b965_iftrue;
     MUX_uxn_c_l311_c44_b965_iffalse <= VAR_MUX_uxn_c_l311_c44_b965_iffalse;
     -- Outputs
     VAR_MUX_uxn_c_l311_c44_b965_return_output := MUX_uxn_c_l311_c44_b965_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_c_l317_c9_9a0e] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_return_output;

     -- Submodule level 2
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_c_l317_c9_9a0e_return_output;
     VAR_MUX_uxn_c_l311_c16_5d3e_iffalse := VAR_MUX_uxn_c_l311_c44_b965_return_output;
     -- MUX[uxn_c_l311_c16_5d3e] LATENCY=0
     -- Inputs
     MUX_uxn_c_l311_c16_5d3e_cond <= VAR_MUX_uxn_c_l311_c16_5d3e_cond;
     MUX_uxn_c_l311_c16_5d3e_iftrue <= VAR_MUX_uxn_c_l311_c16_5d3e_iftrue;
     MUX_uxn_c_l311_c16_5d3e_iffalse <= VAR_MUX_uxn_c_l311_c16_5d3e_iffalse;
     -- Outputs
     VAR_MUX_uxn_c_l311_c16_5d3e_return_output := MUX_uxn_c_l311_c16_5d3e_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_c_l317_c1_20da] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_return_output;

     -- Submodule level 3
     VAR_BIN_OP_EQ_uxn_c_l312_c16_4c21_left := VAR_MUX_uxn_c_l311_c16_5d3e_return_output;
     VAR_boot_check_MUX_uxn_c_l302_c2_9cba_iftrue := VAR_MUX_uxn_c_l311_c16_5d3e_return_output;
     VAR_step_cpu_uxn_c_l318_c21_a9b6_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_c_l317_c1_20da_return_output;
     -- BIN_OP_EQ[uxn_c_l312_c16_4c21] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_c_l312_c16_4c21_left <= VAR_BIN_OP_EQ_uxn_c_l312_c16_4c21_left;
     BIN_OP_EQ_uxn_c_l312_c16_4c21_right <= VAR_BIN_OP_EQ_uxn_c_l312_c16_4c21_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_c_l312_c16_4c21_return_output := BIN_OP_EQ_uxn_c_l312_c16_4c21_return_output;

     -- step_cpu[uxn_c_l318_c21_a9b6] LATENCY=0
     -- Clock enable
     step_cpu_uxn_c_l318_c21_a9b6_CLOCK_ENABLE <= VAR_step_cpu_uxn_c_l318_c21_a9b6_CLOCK_ENABLE;
     -- Inputs
     step_cpu_uxn_c_l318_c21_a9b6_previous_ram_read_value <= VAR_step_cpu_uxn_c_l318_c21_a9b6_previous_ram_read_value;
     step_cpu_uxn_c_l318_c21_a9b6_previous_device_ram_read <= VAR_step_cpu_uxn_c_l318_c21_a9b6_previous_device_ram_read;
     step_cpu_uxn_c_l318_c21_a9b6_use_vector <= VAR_step_cpu_uxn_c_l318_c21_a9b6_use_vector;
     step_cpu_uxn_c_l318_c21_a9b6_vector <= VAR_step_cpu_uxn_c_l318_c21_a9b6_vector;
     -- Outputs
     VAR_step_cpu_uxn_c_l318_c21_a9b6_return_output := step_cpu_uxn_c_l318_c21_a9b6_return_output;

     -- boot_check_MUX[uxn_c_l302_c2_9cba] LATENCY=0
     -- Inputs
     boot_check_MUX_uxn_c_l302_c2_9cba_cond <= VAR_boot_check_MUX_uxn_c_l302_c2_9cba_cond;
     boot_check_MUX_uxn_c_l302_c2_9cba_iftrue <= VAR_boot_check_MUX_uxn_c_l302_c2_9cba_iftrue;
     boot_check_MUX_uxn_c_l302_c2_9cba_iffalse <= VAR_boot_check_MUX_uxn_c_l302_c2_9cba_iffalse;
     -- Outputs
     VAR_boot_check_MUX_uxn_c_l302_c2_9cba_return_output := boot_check_MUX_uxn_c_l302_c2_9cba_return_output;

     -- Submodule level 4
     VAR_MUX_uxn_c_l312_c16_1944_cond := VAR_BIN_OP_EQ_uxn_c_l312_c16_4c21_return_output;
     REG_VAR_boot_check := VAR_boot_check_MUX_uxn_c_l302_c2_9cba_return_output;
     VAR_cpu_step_result_MUX_uxn_c_l317_c9_9a0e_iftrue := VAR_step_cpu_uxn_c_l318_c21_a9b6_return_output;
     -- CONST_REF_RD_uint1_t_cpu_step_result_t_vram_write_layer_d41d[uxn_c_l325_c22_9ead] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_cpu_step_result_t_vram_write_layer_d41d_uxn_c_l325_c22_9ead_return_output := VAR_step_cpu_uxn_c_l318_c21_a9b6_return_output.vram_write_layer;

     -- CONST_REF_RD_uint1_t_cpu_step_result_t_is_ram_write_d41d[uxn_c_l319_c18_e6d8] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_cpu_step_result_t_is_ram_write_d41d_uxn_c_l319_c18_e6d8_return_output := VAR_step_cpu_uxn_c_l318_c21_a9b6_return_output.is_ram_write;

     -- CONST_REF_RD_uint8_t_cpu_step_result_t_device_ram_address_d41d[uxn_c_l321_c24_5ea8] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_cpu_step_result_t_device_ram_address_d41d_uxn_c_l321_c24_5ea8_return_output := VAR_step_cpu_uxn_c_l318_c21_a9b6_return_output.device_ram_address;

     -- CONST_REF_RD_uint1_t_cpu_step_result_t_is_device_ram_write_d41d[uxn_c_l322_c25_df61] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_cpu_step_result_t_is_device_ram_write_d41d_uxn_c_l322_c25_df61_return_output := VAR_step_cpu_uxn_c_l318_c21_a9b6_return_output.is_device_ram_write;

     -- MUX[uxn_c_l312_c16_1944] LATENCY=0
     -- Inputs
     MUX_uxn_c_l312_c16_1944_cond <= VAR_MUX_uxn_c_l312_c16_1944_cond;
     MUX_uxn_c_l312_c16_1944_iftrue <= VAR_MUX_uxn_c_l312_c16_1944_iftrue;
     MUX_uxn_c_l312_c16_1944_iffalse <= VAR_MUX_uxn_c_l312_c16_1944_iffalse;
     -- Outputs
     VAR_MUX_uxn_c_l312_c16_1944_return_output := MUX_uxn_c_l312_c16_1944_return_output;

     -- CONST_REF_RD_uint1_t_cpu_step_result_t_is_vram_write_d41d[uxn_c_l324_c19_bd0b] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_cpu_step_result_t_is_vram_write_d41d_uxn_c_l324_c19_bd0b_return_output := VAR_step_cpu_uxn_c_l318_c21_a9b6_return_output.is_vram_write;

     -- CONST_REF_RD_uint8_t_cpu_step_result_t_u8_value_d41d_uxn_c_l323_l326_DUPLICATE_30f9 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_cpu_step_result_t_u8_value_d41d_uxn_c_l323_l326_DUPLICATE_30f9_return_output := VAR_step_cpu_uxn_c_l318_c21_a9b6_return_output.u8_value;

     -- CONST_REF_RD_uint16_t_cpu_step_result_t_u16_addr_d41d[uxn_c_l320_c14_8d49] LATENCY=0
     VAR_CONST_REF_RD_uint16_t_cpu_step_result_t_u16_addr_d41d_uxn_c_l320_c14_8d49_return_output := VAR_step_cpu_uxn_c_l318_c21_a9b6_return_output.u16_addr;

     -- cpu_step_result_MUX[uxn_c_l317_c9_9a0e] LATENCY=0
     -- Inputs
     cpu_step_result_MUX_uxn_c_l317_c9_9a0e_cond <= VAR_cpu_step_result_MUX_uxn_c_l317_c9_9a0e_cond;
     cpu_step_result_MUX_uxn_c_l317_c9_9a0e_iftrue <= VAR_cpu_step_result_MUX_uxn_c_l317_c9_9a0e_iftrue;
     cpu_step_result_MUX_uxn_c_l317_c9_9a0e_iffalse <= VAR_cpu_step_result_MUX_uxn_c_l317_c9_9a0e_iffalse;
     -- Outputs
     VAR_cpu_step_result_MUX_uxn_c_l317_c9_9a0e_return_output := cpu_step_result_MUX_uxn_c_l317_c9_9a0e_return_output;

     -- Submodule level 5
     VAR_u16_addr_MUX_uxn_c_l317_c9_9a0e_iftrue := VAR_CONST_REF_RD_uint16_t_cpu_step_result_t_u16_addr_d41d_uxn_c_l320_c14_8d49_return_output;
     VAR_is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_iftrue := VAR_CONST_REF_RD_uint1_t_cpu_step_result_t_is_device_ram_write_d41d_uxn_c_l322_c25_df61_return_output;
     VAR_is_ram_write_MUX_uxn_c_l317_c9_9a0e_iftrue := VAR_CONST_REF_RD_uint1_t_cpu_step_result_t_is_ram_write_d41d_uxn_c_l319_c18_e6d8_return_output;
     VAR_is_vram_write_MUX_uxn_c_l317_c9_9a0e_iftrue := VAR_CONST_REF_RD_uint1_t_cpu_step_result_t_is_vram_write_d41d_uxn_c_l324_c19_bd0b_return_output;
     VAR_vram_write_layer_MUX_uxn_c_l317_c9_9a0e_iftrue := VAR_CONST_REF_RD_uint1_t_cpu_step_result_t_vram_write_layer_d41d_uxn_c_l325_c22_9ead_return_output;
     VAR_device_ram_address_MUX_uxn_c_l317_c9_9a0e_iftrue := VAR_CONST_REF_RD_uint8_t_cpu_step_result_t_device_ram_address_d41d_uxn_c_l321_c24_5ea8_return_output;
     VAR_ram_write_value_MUX_uxn_c_l317_c9_9a0e_iftrue := VAR_CONST_REF_RD_uint8_t_cpu_step_result_t_u8_value_d41d_uxn_c_l323_l326_DUPLICATE_30f9_return_output;
     VAR_vram_value_MUX_uxn_c_l317_c9_9a0e_iftrue := VAR_CONST_REF_RD_uint8_t_cpu_step_result_t_u8_value_d41d_uxn_c_l323_l326_DUPLICATE_30f9_return_output;
     VAR_BIN_OP_OR_uint1_t_uint1_t_uxn_c_l313_l314_DUPLICATE_e2dd_right := VAR_MUX_uxn_c_l312_c16_1944_return_output;
     VAR_MUX_uxn_c_l315_c21_ddb1_cond := VAR_MUX_uxn_c_l312_c16_1944_return_output;
     VAR_is_booted_MUX_uxn_c_l302_c2_9cba_iftrue := VAR_MUX_uxn_c_l312_c16_1944_return_output;
     VAR_cpu_step_result_MUX_uxn_c_l302_c2_9cba_iffalse := VAR_cpu_step_result_MUX_uxn_c_l317_c9_9a0e_return_output;
     -- is_ram_write_MUX[uxn_c_l317_c9_9a0e] LATENCY=0
     -- Inputs
     is_ram_write_MUX_uxn_c_l317_c9_9a0e_cond <= VAR_is_ram_write_MUX_uxn_c_l317_c9_9a0e_cond;
     is_ram_write_MUX_uxn_c_l317_c9_9a0e_iftrue <= VAR_is_ram_write_MUX_uxn_c_l317_c9_9a0e_iftrue;
     is_ram_write_MUX_uxn_c_l317_c9_9a0e_iffalse <= VAR_is_ram_write_MUX_uxn_c_l317_c9_9a0e_iffalse;
     -- Outputs
     VAR_is_ram_write_MUX_uxn_c_l317_c9_9a0e_return_output := is_ram_write_MUX_uxn_c_l317_c9_9a0e_return_output;

     -- u16_addr_MUX[uxn_c_l317_c9_9a0e] LATENCY=0
     -- Inputs
     u16_addr_MUX_uxn_c_l317_c9_9a0e_cond <= VAR_u16_addr_MUX_uxn_c_l317_c9_9a0e_cond;
     u16_addr_MUX_uxn_c_l317_c9_9a0e_iftrue <= VAR_u16_addr_MUX_uxn_c_l317_c9_9a0e_iftrue;
     u16_addr_MUX_uxn_c_l317_c9_9a0e_iffalse <= VAR_u16_addr_MUX_uxn_c_l317_c9_9a0e_iffalse;
     -- Outputs
     VAR_u16_addr_MUX_uxn_c_l317_c9_9a0e_return_output := u16_addr_MUX_uxn_c_l317_c9_9a0e_return_output;

     -- vram_value_MUX[uxn_c_l317_c9_9a0e] LATENCY=0
     -- Inputs
     vram_value_MUX_uxn_c_l317_c9_9a0e_cond <= VAR_vram_value_MUX_uxn_c_l317_c9_9a0e_cond;
     vram_value_MUX_uxn_c_l317_c9_9a0e_iftrue <= VAR_vram_value_MUX_uxn_c_l317_c9_9a0e_iftrue;
     vram_value_MUX_uxn_c_l317_c9_9a0e_iffalse <= VAR_vram_value_MUX_uxn_c_l317_c9_9a0e_iffalse;
     -- Outputs
     VAR_vram_value_MUX_uxn_c_l317_c9_9a0e_return_output := vram_value_MUX_uxn_c_l317_c9_9a0e_return_output;

     -- is_device_ram_write_MUX[uxn_c_l317_c9_9a0e] LATENCY=0
     -- Inputs
     is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_cond <= VAR_is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_cond;
     is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_iftrue <= VAR_is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_iftrue;
     is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_iffalse <= VAR_is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_iffalse;
     -- Outputs
     VAR_is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_return_output := is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_return_output;

     -- BIN_OP_OR_uint1_t_uint1_t_uxn_c_l313_l314_DUPLICATE_e2dd LATENCY=0
     -- Inputs
     BIN_OP_OR_uint1_t_uint1_t_uxn_c_l313_l314_DUPLICATE_e2dd_left <= VAR_BIN_OP_OR_uint1_t_uint1_t_uxn_c_l313_l314_DUPLICATE_e2dd_left;
     BIN_OP_OR_uint1_t_uint1_t_uxn_c_l313_l314_DUPLICATE_e2dd_right <= VAR_BIN_OP_OR_uint1_t_uint1_t_uxn_c_l313_l314_DUPLICATE_e2dd_right;
     -- Outputs
     VAR_BIN_OP_OR_uint1_t_uint1_t_uxn_c_l313_l314_DUPLICATE_e2dd_return_output := BIN_OP_OR_uint1_t_uint1_t_uxn_c_l313_l314_DUPLICATE_e2dd_return_output;

     -- is_vram_write_MUX[uxn_c_l317_c9_9a0e] LATENCY=0
     -- Inputs
     is_vram_write_MUX_uxn_c_l317_c9_9a0e_cond <= VAR_is_vram_write_MUX_uxn_c_l317_c9_9a0e_cond;
     is_vram_write_MUX_uxn_c_l317_c9_9a0e_iftrue <= VAR_is_vram_write_MUX_uxn_c_l317_c9_9a0e_iftrue;
     is_vram_write_MUX_uxn_c_l317_c9_9a0e_iffalse <= VAR_is_vram_write_MUX_uxn_c_l317_c9_9a0e_iffalse;
     -- Outputs
     VAR_is_vram_write_MUX_uxn_c_l317_c9_9a0e_return_output := is_vram_write_MUX_uxn_c_l317_c9_9a0e_return_output;

     -- device_ram_address_MUX[uxn_c_l317_c9_9a0e] LATENCY=0
     -- Inputs
     device_ram_address_MUX_uxn_c_l317_c9_9a0e_cond <= VAR_device_ram_address_MUX_uxn_c_l317_c9_9a0e_cond;
     device_ram_address_MUX_uxn_c_l317_c9_9a0e_iftrue <= VAR_device_ram_address_MUX_uxn_c_l317_c9_9a0e_iftrue;
     device_ram_address_MUX_uxn_c_l317_c9_9a0e_iffalse <= VAR_device_ram_address_MUX_uxn_c_l317_c9_9a0e_iffalse;
     -- Outputs
     VAR_device_ram_address_MUX_uxn_c_l317_c9_9a0e_return_output := device_ram_address_MUX_uxn_c_l317_c9_9a0e_return_output;

     -- MUX[uxn_c_l315_c21_ddb1] LATENCY=0
     -- Inputs
     MUX_uxn_c_l315_c21_ddb1_cond <= VAR_MUX_uxn_c_l315_c21_ddb1_cond;
     MUX_uxn_c_l315_c21_ddb1_iftrue <= VAR_MUX_uxn_c_l315_c21_ddb1_iftrue;
     MUX_uxn_c_l315_c21_ddb1_iffalse <= VAR_MUX_uxn_c_l315_c21_ddb1_iffalse;
     -- Outputs
     VAR_MUX_uxn_c_l315_c21_ddb1_return_output := MUX_uxn_c_l315_c21_ddb1_return_output;

     -- ram_write_value_MUX[uxn_c_l317_c9_9a0e] LATENCY=0
     -- Inputs
     ram_write_value_MUX_uxn_c_l317_c9_9a0e_cond <= VAR_ram_write_value_MUX_uxn_c_l317_c9_9a0e_cond;
     ram_write_value_MUX_uxn_c_l317_c9_9a0e_iftrue <= VAR_ram_write_value_MUX_uxn_c_l317_c9_9a0e_iftrue;
     ram_write_value_MUX_uxn_c_l317_c9_9a0e_iffalse <= VAR_ram_write_value_MUX_uxn_c_l317_c9_9a0e_iffalse;
     -- Outputs
     VAR_ram_write_value_MUX_uxn_c_l317_c9_9a0e_return_output := ram_write_value_MUX_uxn_c_l317_c9_9a0e_return_output;

     -- cpu_step_result_MUX[uxn_c_l302_c2_9cba] LATENCY=0
     -- Inputs
     cpu_step_result_MUX_uxn_c_l302_c2_9cba_cond <= VAR_cpu_step_result_MUX_uxn_c_l302_c2_9cba_cond;
     cpu_step_result_MUX_uxn_c_l302_c2_9cba_iftrue <= VAR_cpu_step_result_MUX_uxn_c_l302_c2_9cba_iftrue;
     cpu_step_result_MUX_uxn_c_l302_c2_9cba_iffalse <= VAR_cpu_step_result_MUX_uxn_c_l302_c2_9cba_iffalse;
     -- Outputs
     VAR_cpu_step_result_MUX_uxn_c_l302_c2_9cba_return_output := cpu_step_result_MUX_uxn_c_l302_c2_9cba_return_output;

     -- vram_write_layer_MUX[uxn_c_l317_c9_9a0e] LATENCY=0
     -- Inputs
     vram_write_layer_MUX_uxn_c_l317_c9_9a0e_cond <= VAR_vram_write_layer_MUX_uxn_c_l317_c9_9a0e_cond;
     vram_write_layer_MUX_uxn_c_l317_c9_9a0e_iftrue <= VAR_vram_write_layer_MUX_uxn_c_l317_c9_9a0e_iftrue;
     vram_write_layer_MUX_uxn_c_l317_c9_9a0e_iffalse <= VAR_vram_write_layer_MUX_uxn_c_l317_c9_9a0e_iffalse;
     -- Outputs
     VAR_vram_write_layer_MUX_uxn_c_l317_c9_9a0e_return_output := vram_write_layer_MUX_uxn_c_l317_c9_9a0e_return_output;

     -- is_booted_MUX[uxn_c_l302_c2_9cba] LATENCY=0
     -- Inputs
     is_booted_MUX_uxn_c_l302_c2_9cba_cond <= VAR_is_booted_MUX_uxn_c_l302_c2_9cba_cond;
     is_booted_MUX_uxn_c_l302_c2_9cba_iftrue <= VAR_is_booted_MUX_uxn_c_l302_c2_9cba_iftrue;
     is_booted_MUX_uxn_c_l302_c2_9cba_iffalse <= VAR_is_booted_MUX_uxn_c_l302_c2_9cba_iffalse;
     -- Outputs
     VAR_is_booted_MUX_uxn_c_l302_c2_9cba_return_output := is_booted_MUX_uxn_c_l302_c2_9cba_return_output;

     -- Submodule level 6
     VAR_MUX_uxn_c_l314_c16_61c4_cond := VAR_BIN_OP_OR_uint1_t_uint1_t_uxn_c_l313_l314_DUPLICATE_e2dd_return_output;
     VAR_is_ram_write_MUX_uxn_c_l302_c2_9cba_iftrue := VAR_BIN_OP_OR_uint1_t_uint1_t_uxn_c_l313_l314_DUPLICATE_e2dd_return_output;
     VAR_ram_write_value_MUX_uxn_c_l302_c2_9cba_iftrue := VAR_MUX_uxn_c_l315_c21_ddb1_return_output;
     REG_VAR_cpu_step_result := VAR_cpu_step_result_MUX_uxn_c_l302_c2_9cba_return_output;
     VAR_device_ram_address_MUX_uxn_c_l302_c2_9cba_iffalse := VAR_device_ram_address_MUX_uxn_c_l317_c9_9a0e_return_output;
     REG_VAR_is_booted := VAR_is_booted_MUX_uxn_c_l302_c2_9cba_return_output;
     VAR_is_device_ram_write_MUX_uxn_c_l302_c2_9cba_iffalse := VAR_is_device_ram_write_MUX_uxn_c_l317_c9_9a0e_return_output;
     VAR_is_ram_write_MUX_uxn_c_l302_c2_9cba_iffalse := VAR_is_ram_write_MUX_uxn_c_l317_c9_9a0e_return_output;
     VAR_is_vram_write_MUX_uxn_c_l302_c2_9cba_iffalse := VAR_is_vram_write_MUX_uxn_c_l317_c9_9a0e_return_output;
     VAR_ram_write_value_MUX_uxn_c_l302_c2_9cba_iffalse := VAR_ram_write_value_MUX_uxn_c_l317_c9_9a0e_return_output;
     VAR_u16_addr_MUX_uxn_c_l302_c2_9cba_iffalse := VAR_u16_addr_MUX_uxn_c_l317_c9_9a0e_return_output;
     VAR_vram_value_MUX_uxn_c_l302_c2_9cba_iffalse := VAR_vram_value_MUX_uxn_c_l317_c9_9a0e_return_output;
     VAR_vram_write_layer_MUX_uxn_c_l302_c2_9cba_iffalse := VAR_vram_write_layer_MUX_uxn_c_l317_c9_9a0e_return_output;
     -- is_device_ram_write_MUX[uxn_c_l302_c2_9cba] LATENCY=0
     -- Inputs
     is_device_ram_write_MUX_uxn_c_l302_c2_9cba_cond <= VAR_is_device_ram_write_MUX_uxn_c_l302_c2_9cba_cond;
     is_device_ram_write_MUX_uxn_c_l302_c2_9cba_iftrue <= VAR_is_device_ram_write_MUX_uxn_c_l302_c2_9cba_iftrue;
     is_device_ram_write_MUX_uxn_c_l302_c2_9cba_iffalse <= VAR_is_device_ram_write_MUX_uxn_c_l302_c2_9cba_iffalse;
     -- Outputs
     VAR_is_device_ram_write_MUX_uxn_c_l302_c2_9cba_return_output := is_device_ram_write_MUX_uxn_c_l302_c2_9cba_return_output;

     -- is_ram_write_MUX[uxn_c_l302_c2_9cba] LATENCY=0
     -- Inputs
     is_ram_write_MUX_uxn_c_l302_c2_9cba_cond <= VAR_is_ram_write_MUX_uxn_c_l302_c2_9cba_cond;
     is_ram_write_MUX_uxn_c_l302_c2_9cba_iftrue <= VAR_is_ram_write_MUX_uxn_c_l302_c2_9cba_iftrue;
     is_ram_write_MUX_uxn_c_l302_c2_9cba_iffalse <= VAR_is_ram_write_MUX_uxn_c_l302_c2_9cba_iffalse;
     -- Outputs
     VAR_is_ram_write_MUX_uxn_c_l302_c2_9cba_return_output := is_ram_write_MUX_uxn_c_l302_c2_9cba_return_output;

     -- device_ram_address_MUX[uxn_c_l302_c2_9cba] LATENCY=0
     -- Inputs
     device_ram_address_MUX_uxn_c_l302_c2_9cba_cond <= VAR_device_ram_address_MUX_uxn_c_l302_c2_9cba_cond;
     device_ram_address_MUX_uxn_c_l302_c2_9cba_iftrue <= VAR_device_ram_address_MUX_uxn_c_l302_c2_9cba_iftrue;
     device_ram_address_MUX_uxn_c_l302_c2_9cba_iffalse <= VAR_device_ram_address_MUX_uxn_c_l302_c2_9cba_iffalse;
     -- Outputs
     VAR_device_ram_address_MUX_uxn_c_l302_c2_9cba_return_output := device_ram_address_MUX_uxn_c_l302_c2_9cba_return_output;

     -- is_vram_write_MUX[uxn_c_l302_c2_9cba] LATENCY=0
     -- Inputs
     is_vram_write_MUX_uxn_c_l302_c2_9cba_cond <= VAR_is_vram_write_MUX_uxn_c_l302_c2_9cba_cond;
     is_vram_write_MUX_uxn_c_l302_c2_9cba_iftrue <= VAR_is_vram_write_MUX_uxn_c_l302_c2_9cba_iftrue;
     is_vram_write_MUX_uxn_c_l302_c2_9cba_iffalse <= VAR_is_vram_write_MUX_uxn_c_l302_c2_9cba_iffalse;
     -- Outputs
     VAR_is_vram_write_MUX_uxn_c_l302_c2_9cba_return_output := is_vram_write_MUX_uxn_c_l302_c2_9cba_return_output;

     -- vram_value_MUX[uxn_c_l302_c2_9cba] LATENCY=0
     -- Inputs
     vram_value_MUX_uxn_c_l302_c2_9cba_cond <= VAR_vram_value_MUX_uxn_c_l302_c2_9cba_cond;
     vram_value_MUX_uxn_c_l302_c2_9cba_iftrue <= VAR_vram_value_MUX_uxn_c_l302_c2_9cba_iftrue;
     vram_value_MUX_uxn_c_l302_c2_9cba_iffalse <= VAR_vram_value_MUX_uxn_c_l302_c2_9cba_iffalse;
     -- Outputs
     VAR_vram_value_MUX_uxn_c_l302_c2_9cba_return_output := vram_value_MUX_uxn_c_l302_c2_9cba_return_output;

     -- ram_write_value_MUX[uxn_c_l302_c2_9cba] LATENCY=0
     -- Inputs
     ram_write_value_MUX_uxn_c_l302_c2_9cba_cond <= VAR_ram_write_value_MUX_uxn_c_l302_c2_9cba_cond;
     ram_write_value_MUX_uxn_c_l302_c2_9cba_iftrue <= VAR_ram_write_value_MUX_uxn_c_l302_c2_9cba_iftrue;
     ram_write_value_MUX_uxn_c_l302_c2_9cba_iffalse <= VAR_ram_write_value_MUX_uxn_c_l302_c2_9cba_iffalse;
     -- Outputs
     VAR_ram_write_value_MUX_uxn_c_l302_c2_9cba_return_output := ram_write_value_MUX_uxn_c_l302_c2_9cba_return_output;

     -- MUX[uxn_c_l314_c16_61c4] LATENCY=0
     -- Inputs
     MUX_uxn_c_l314_c16_61c4_cond <= VAR_MUX_uxn_c_l314_c16_61c4_cond;
     MUX_uxn_c_l314_c16_61c4_iftrue <= VAR_MUX_uxn_c_l314_c16_61c4_iftrue;
     MUX_uxn_c_l314_c16_61c4_iffalse <= VAR_MUX_uxn_c_l314_c16_61c4_iffalse;
     -- Outputs
     VAR_MUX_uxn_c_l314_c16_61c4_return_output := MUX_uxn_c_l314_c16_61c4_return_output;

     -- vram_write_layer_MUX[uxn_c_l302_c2_9cba] LATENCY=0
     -- Inputs
     vram_write_layer_MUX_uxn_c_l302_c2_9cba_cond <= VAR_vram_write_layer_MUX_uxn_c_l302_c2_9cba_cond;
     vram_write_layer_MUX_uxn_c_l302_c2_9cba_iftrue <= VAR_vram_write_layer_MUX_uxn_c_l302_c2_9cba_iftrue;
     vram_write_layer_MUX_uxn_c_l302_c2_9cba_iffalse <= VAR_vram_write_layer_MUX_uxn_c_l302_c2_9cba_iffalse;
     -- Outputs
     VAR_vram_write_layer_MUX_uxn_c_l302_c2_9cba_return_output := vram_write_layer_MUX_uxn_c_l302_c2_9cba_return_output;

     -- Submodule level 7
     VAR_BIN_OP_PLUS_uxn_c_l314_c3_4639_right := VAR_MUX_uxn_c_l314_c16_61c4_return_output;
     REG_VAR_device_ram_address := VAR_device_ram_address_MUX_uxn_c_l302_c2_9cba_return_output;
     VAR_device_ram_update_uxn_c_l335_c26_db12_device_address := VAR_device_ram_address_MUX_uxn_c_l302_c2_9cba_return_output;
     VAR_palette_snoop_uxn_c_l343_c20_f328_device_ram_address := VAR_device_ram_address_MUX_uxn_c_l302_c2_9cba_return_output;
     VAR_vector_snoop_uxn_c_l344_c18_80ab_device_ram_address := VAR_device_ram_address_MUX_uxn_c_l302_c2_9cba_return_output;
     VAR_device_ram_update_uxn_c_l335_c26_db12_write_enable := VAR_is_device_ram_write_MUX_uxn_c_l302_c2_9cba_return_output;
     REG_VAR_is_device_ram_write := VAR_is_device_ram_write_MUX_uxn_c_l302_c2_9cba_return_output;
     VAR_palette_snoop_uxn_c_l343_c20_f328_is_device_ram_write := VAR_is_device_ram_write_MUX_uxn_c_l302_c2_9cba_return_output;
     VAR_vector_snoop_uxn_c_l344_c18_80ab_is_device_ram_write := VAR_is_device_ram_write_MUX_uxn_c_l302_c2_9cba_return_output;
     REG_VAR_is_ram_write := VAR_is_ram_write_MUX_uxn_c_l302_c2_9cba_return_output;
     VAR_main_ram_update_uxn_c_l329_c19_6697_write_enable := VAR_is_ram_write_MUX_uxn_c_l302_c2_9cba_return_output;
     REG_VAR_is_vram_write := VAR_is_vram_write_MUX_uxn_c_l302_c2_9cba_return_output;
     VAR_step_gpu_uxn_c_l341_c20_9854_is_vram_write := VAR_is_vram_write_MUX_uxn_c_l302_c2_9cba_return_output;
     VAR_device_ram_update_uxn_c_l335_c26_db12_value := VAR_ram_write_value_MUX_uxn_c_l302_c2_9cba_return_output;
     VAR_main_ram_update_uxn_c_l329_c19_6697_value := VAR_ram_write_value_MUX_uxn_c_l302_c2_9cba_return_output;
     VAR_palette_snoop_uxn_c_l343_c20_f328_device_ram_value := VAR_ram_write_value_MUX_uxn_c_l302_c2_9cba_return_output;
     REG_VAR_ram_write_value := VAR_ram_write_value_MUX_uxn_c_l302_c2_9cba_return_output;
     VAR_vector_snoop_uxn_c_l344_c18_80ab_device_ram_value := VAR_ram_write_value_MUX_uxn_c_l302_c2_9cba_return_output;
     VAR_step_gpu_uxn_c_l341_c20_9854_vram_value := VAR_vram_value_MUX_uxn_c_l302_c2_9cba_return_output;
     REG_VAR_vram_value := VAR_vram_value_MUX_uxn_c_l302_c2_9cba_return_output;
     VAR_step_gpu_uxn_c_l341_c20_9854_vram_write_layer := VAR_vram_write_layer_MUX_uxn_c_l302_c2_9cba_return_output;
     REG_VAR_vram_write_layer := VAR_vram_write_layer_MUX_uxn_c_l302_c2_9cba_return_output;
     -- BIN_OP_PLUS[uxn_c_l314_c3_4639] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_c_l314_c3_4639_left <= VAR_BIN_OP_PLUS_uxn_c_l314_c3_4639_left;
     BIN_OP_PLUS_uxn_c_l314_c3_4639_right <= VAR_BIN_OP_PLUS_uxn_c_l314_c3_4639_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_c_l314_c3_4639_return_output := BIN_OP_PLUS_uxn_c_l314_c3_4639_return_output;

     -- vector_snoop[uxn_c_l344_c18_80ab] LATENCY=0
     -- Clock enable
     vector_snoop_uxn_c_l344_c18_80ab_CLOCK_ENABLE <= VAR_vector_snoop_uxn_c_l344_c18_80ab_CLOCK_ENABLE;
     -- Inputs
     vector_snoop_uxn_c_l344_c18_80ab_device_ram_address <= VAR_vector_snoop_uxn_c_l344_c18_80ab_device_ram_address;
     vector_snoop_uxn_c_l344_c18_80ab_device_ram_value <= VAR_vector_snoop_uxn_c_l344_c18_80ab_device_ram_value;
     vector_snoop_uxn_c_l344_c18_80ab_is_device_ram_write <= VAR_vector_snoop_uxn_c_l344_c18_80ab_is_device_ram_write;
     -- Outputs
     VAR_vector_snoop_uxn_c_l344_c18_80ab_return_output := vector_snoop_uxn_c_l344_c18_80ab_return_output;

     -- device_ram_update[uxn_c_l335_c26_db12] LATENCY=0
     -- Clock enable
     device_ram_update_uxn_c_l335_c26_db12_CLOCK_ENABLE <= VAR_device_ram_update_uxn_c_l335_c26_db12_CLOCK_ENABLE;
     -- Inputs
     device_ram_update_uxn_c_l335_c26_db12_device_address <= VAR_device_ram_update_uxn_c_l335_c26_db12_device_address;
     device_ram_update_uxn_c_l335_c26_db12_value <= VAR_device_ram_update_uxn_c_l335_c26_db12_value;
     device_ram_update_uxn_c_l335_c26_db12_write_enable <= VAR_device_ram_update_uxn_c_l335_c26_db12_write_enable;
     -- Outputs
     VAR_device_ram_update_uxn_c_l335_c26_db12_return_output := device_ram_update_uxn_c_l335_c26_db12_return_output;

     -- Submodule level 8
     VAR_u16_addr_uxn_c_l314_c3_4336 := resize(VAR_BIN_OP_PLUS_uxn_c_l314_c3_4639_return_output, 16);
     REG_VAR_device_ram_read_value := VAR_device_ram_update_uxn_c_l335_c26_db12_return_output;
     REG_VAR_screen_vector := VAR_vector_snoop_uxn_c_l344_c18_80ab_return_output;
     VAR_u16_addr_MUX_uxn_c_l302_c2_9cba_iftrue := VAR_u16_addr_uxn_c_l314_c3_4336;
     -- u16_addr_MUX[uxn_c_l302_c2_9cba] LATENCY=0
     -- Inputs
     u16_addr_MUX_uxn_c_l302_c2_9cba_cond <= VAR_u16_addr_MUX_uxn_c_l302_c2_9cba_cond;
     u16_addr_MUX_uxn_c_l302_c2_9cba_iftrue <= VAR_u16_addr_MUX_uxn_c_l302_c2_9cba_iftrue;
     u16_addr_MUX_uxn_c_l302_c2_9cba_iffalse <= VAR_u16_addr_MUX_uxn_c_l302_c2_9cba_iffalse;
     -- Outputs
     VAR_u16_addr_MUX_uxn_c_l302_c2_9cba_return_output := u16_addr_MUX_uxn_c_l302_c2_9cba_return_output;

     -- Submodule level 9
     VAR_main_ram_update_uxn_c_l329_c19_6697_ram_address := VAR_u16_addr_MUX_uxn_c_l302_c2_9cba_return_output;
     VAR_step_gpu_uxn_c_l341_c20_9854_vram_address := VAR_u16_addr_MUX_uxn_c_l302_c2_9cba_return_output;
     REG_VAR_u16_addr := VAR_u16_addr_MUX_uxn_c_l302_c2_9cba_return_output;
     -- main_ram_update[uxn_c_l329_c19_6697] LATENCY=0
     -- Clock enable
     main_ram_update_uxn_c_l329_c19_6697_CLOCK_ENABLE <= VAR_main_ram_update_uxn_c_l329_c19_6697_CLOCK_ENABLE;
     -- Inputs
     main_ram_update_uxn_c_l329_c19_6697_ram_address <= VAR_main_ram_update_uxn_c_l329_c19_6697_ram_address;
     main_ram_update_uxn_c_l329_c19_6697_value <= VAR_main_ram_update_uxn_c_l329_c19_6697_value;
     main_ram_update_uxn_c_l329_c19_6697_write_enable <= VAR_main_ram_update_uxn_c_l329_c19_6697_write_enable;
     -- Outputs
     VAR_main_ram_update_uxn_c_l329_c19_6697_return_output := main_ram_update_uxn_c_l329_c19_6697_return_output;

     -- step_gpu[uxn_c_l341_c20_9854] LATENCY=0
     -- Clock enable
     step_gpu_uxn_c_l341_c20_9854_CLOCK_ENABLE <= VAR_step_gpu_uxn_c_l341_c20_9854_CLOCK_ENABLE;
     -- Inputs
     step_gpu_uxn_c_l341_c20_9854_is_active_drawing_area <= VAR_step_gpu_uxn_c_l341_c20_9854_is_active_drawing_area;
     step_gpu_uxn_c_l341_c20_9854_is_vram_write <= VAR_step_gpu_uxn_c_l341_c20_9854_is_vram_write;
     step_gpu_uxn_c_l341_c20_9854_vram_write_layer <= VAR_step_gpu_uxn_c_l341_c20_9854_vram_write_layer;
     step_gpu_uxn_c_l341_c20_9854_vram_address <= VAR_step_gpu_uxn_c_l341_c20_9854_vram_address;
     step_gpu_uxn_c_l341_c20_9854_vram_value <= VAR_step_gpu_uxn_c_l341_c20_9854_vram_value;
     -- Outputs
     VAR_step_gpu_uxn_c_l341_c20_9854_return_output := step_gpu_uxn_c_l341_c20_9854_return_output;

     -- Submodule level 10
     REG_VAR_ram_read_value := VAR_main_ram_update_uxn_c_l329_c19_6697_return_output;
     REG_VAR_gpu_step_result := VAR_step_gpu_uxn_c_l341_c20_9854_return_output;
     -- CONST_REF_RD_uint2_t_gpu_step_result_t_color_d41d[uxn_c_l343_c92_ec5c] LATENCY=0
     VAR_CONST_REF_RD_uint2_t_gpu_step_result_t_color_d41d_uxn_c_l343_c92_ec5c_return_output := VAR_step_gpu_uxn_c_l341_c20_9854_return_output.color;

     -- CONST_REF_RD_uint1_t_gpu_step_result_t_is_active_fill_d41d[uxn_c_l342_c19_b60d] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_gpu_step_result_t_is_active_fill_d41d_uxn_c_l342_c19_b60d_return_output := VAR_step_gpu_uxn_c_l341_c20_9854_return_output.is_active_fill;

     -- Submodule level 11
     REG_VAR_is_active_fill := VAR_CONST_REF_RD_uint1_t_gpu_step_result_t_is_active_fill_d41d_uxn_c_l342_c19_b60d_return_output;
     VAR_palette_snoop_uxn_c_l343_c20_f328_gpu_step_color := VAR_CONST_REF_RD_uint2_t_gpu_step_result_t_color_d41d_uxn_c_l343_c92_ec5c_return_output;
     -- palette_snoop[uxn_c_l343_c20_f328] LATENCY=0
     -- Clock enable
     palette_snoop_uxn_c_l343_c20_f328_CLOCK_ENABLE <= VAR_palette_snoop_uxn_c_l343_c20_f328_CLOCK_ENABLE;
     -- Inputs
     palette_snoop_uxn_c_l343_c20_f328_device_ram_address <= VAR_palette_snoop_uxn_c_l343_c20_f328_device_ram_address;
     palette_snoop_uxn_c_l343_c20_f328_device_ram_value <= VAR_palette_snoop_uxn_c_l343_c20_f328_device_ram_value;
     palette_snoop_uxn_c_l343_c20_f328_is_device_ram_write <= VAR_palette_snoop_uxn_c_l343_c20_f328_is_device_ram_write;
     palette_snoop_uxn_c_l343_c20_f328_gpu_step_color <= VAR_palette_snoop_uxn_c_l343_c20_f328_gpu_step_color;
     -- Outputs
     VAR_palette_snoop_uxn_c_l343_c20_f328_return_output := palette_snoop_uxn_c_l343_c20_f328_return_output;

     -- Submodule level 12
     VAR_return_output := VAR_palette_snoop_uxn_c_l343_c20_f328_return_output;
     REG_VAR_uxn_eval_result := VAR_palette_snoop_uxn_c_l343_c20_f328_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_boot_check <= REG_VAR_boot_check;
REG_COMB_uxn_eval_result <= REG_VAR_uxn_eval_result;
REG_COMB_is_booted <= REG_VAR_is_booted;
REG_COMB_gpu_step_result <= REG_VAR_gpu_step_result;
REG_COMB_cpu_step_result <= REG_VAR_cpu_step_result;
REG_COMB_is_active_fill <= REG_VAR_is_active_fill;
REG_COMB_is_ram_write <= REG_VAR_is_ram_write;
REG_COMB_u16_addr <= REG_VAR_u16_addr;
REG_COMB_screen_vector <= REG_VAR_screen_vector;
REG_COMB_ram_write_value <= REG_VAR_ram_write_value;
REG_COMB_ram_read_value <= REG_VAR_ram_read_value;
REG_COMB_device_ram_address <= REG_VAR_device_ram_address;
REG_COMB_device_ram_read_value <= REG_VAR_device_ram_read_value;
REG_COMB_is_device_ram_write <= REG_VAR_is_device_ram_write;
REG_COMB_is_vram_write <= REG_VAR_is_vram_write;
REG_COMB_vram_write_layer <= REG_VAR_vram_write_layer;
REG_COMB_vram_value <= REG_VAR_vram_value;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     boot_check <= REG_COMB_boot_check;
     uxn_eval_result <= REG_COMB_uxn_eval_result;
     is_booted <= REG_COMB_is_booted;
     gpu_step_result <= REG_COMB_gpu_step_result;
     cpu_step_result <= REG_COMB_cpu_step_result;
     is_active_fill <= REG_COMB_is_active_fill;
     is_ram_write <= REG_COMB_is_ram_write;
     u16_addr <= REG_COMB_u16_addr;
     screen_vector <= REG_COMB_screen_vector;
     ram_write_value <= REG_COMB_ram_write_value;
     ram_read_value <= REG_COMB_ram_read_value;
     device_ram_address <= REG_COMB_device_ram_address;
     device_ram_read_value <= REG_COMB_device_ram_read_value;
     is_device_ram_write <= REG_COMB_is_device_ram_write;
     is_vram_write <= REG_COMB_is_vram_write;
     vram_write_layer <= REG_COMB_vram_write_layer;
     vram_value <= REG_COMB_vram_value;
 end if;
 end if;
end process;

end arch;
