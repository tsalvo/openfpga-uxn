-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 36
entity nip2_0CLK_1a2ef46d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end nip2_0CLK_1a2ef46d;
architecture arch of nip2_0CLK_1a2ef46d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2174_c6_8acd]
signal BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2174_c2_0f61]
signal t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2174_c2_0f61]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output : signed(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2174_c2_0f61]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2174_c2_0f61]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2174_c2_0f61]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2174_c2_0f61]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output : unsigned(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2174_c2_0f61]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2174_c2_0f61]
signal result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2174_c2_0f61]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2174_c2_0f61]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2174_c2_0f61]
signal t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2187_c11_e301]
signal BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2187_c7_85f5]
signal t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2187_c7_85f5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2187_c7_85f5]
signal result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2187_c7_85f5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2187_c7_85f5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2187_c7_85f5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output : unsigned(3 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2187_c7_85f5]
signal t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2190_c11_25ae]
signal BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2190_c7_8b8e]
signal t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2190_c7_8b8e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2190_c7_8b8e]
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2190_c7_8b8e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2190_c7_8b8e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2190_c7_8b8e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output : unsigned(3 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2190_c7_8b8e]
signal t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2192_c30_e0af]
signal sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2197_c11_5956]
signal BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2197_c7_47bd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2197_c7_47bd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2197_c7_47bd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2197_c7_47bd]
signal result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output : unsigned(7 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2197_c7_47bd]
signal t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_ee25( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.is_vram_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd
BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_left,
BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_right,
BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61
t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_cond,
t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue,
t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse,
t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61
result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61
result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61
result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61
result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61
result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_cond,
result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61
result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61
result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61
t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_cond,
t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue,
t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse,
t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301
BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_left,
BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_right,
BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5
t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_cond,
t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue,
t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse,
t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_cond,
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5
t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_cond,
t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue,
t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse,
t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae
BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_left,
BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_right,
BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e
t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond,
t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue,
t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse,
t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond,
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e
t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond,
t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue,
t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse,
t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af
sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_ins,
sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_x,
sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_y,
sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956
BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956_left,
BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956_right,
BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_cond,
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd
t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_cond,
t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue,
t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse,
t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_return_output,
 t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output,
 t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_return_output,
 t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output,
 t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_return_output,
 t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output,
 t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output,
 sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output,
 t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_return_output : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2179_c3_83e2 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2174_c2_0f61_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2184_c3_cf5e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2174_c2_0f61_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2174_c2_0f61_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2174_c2_0f61_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_return_output : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2188_c3_0f8a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_return_output : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2194_c3_b85b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2199_c3_cead : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2200_c3_cb79 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2197_c7_47bd_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2187_l2174_l2197_DUPLICATE_e1af_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2187_l2197_DUPLICATE_9216_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_2cd6_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2187_l2190_l2197_DUPLICATE_ca71_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ee25_uxn_opcodes_h_l2205_l2170_DUPLICATE_7b84_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2179_c3_83e2 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2179_c3_83e2;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2199_c3_cead := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2199_c3_cead;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_y := resize(to_signed(-2, 3), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2184_c3_cf5e := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2184_c3_cf5e;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2200_c3_cb79 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2200_c3_cb79;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2194_c3_b85b := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2194_c3_b85b;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_right := to_unsigned(2, 2);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2188_c3_0f8a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2188_c3_0f8a;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_right := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue := VAR_previous_stack_read;
     VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse := t16_high;
     VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse := t16_low;
     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2197_c7_47bd] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2197_c7_47bd_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2187_l2197_DUPLICATE_9216 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2187_l2197_DUPLICATE_9216_return_output := result.sp_relative_shift;

     -- sp_relative_shift[uxn_opcodes_h_l2192_c30_e0af] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_ins;
     sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_x;
     sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_return_output := sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2187_l2190_l2197_DUPLICATE_ca71 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2187_l2190_l2197_DUPLICATE_ca71_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2190_c11_25ae] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_left;
     BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_return_output := BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_2cd6 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_2cd6_return_output := result.is_stack_write;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2174_c2_0f61] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2174_c2_0f61_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2174_c6_8acd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_left;
     BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_return_output := BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2197_c11_5956] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956_left;
     BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956_return_output := BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2187_c11_e301] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_left;
     BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_return_output := BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2174_c2_0f61] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2174_c2_0f61_return_output := result.is_stack_index_flipped;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2174_c2_0f61] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2174_c2_0f61_return_output := result.is_pc_updated;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2174_c2_0f61] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2174_c2_0f61_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2187_l2174_l2197_DUPLICATE_e1af LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2187_l2174_l2197_DUPLICATE_e1af_return_output := result.u8_value;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_8acd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_e301_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_25ae_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_5956_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2187_l2197_DUPLICATE_9216_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2187_l2197_DUPLICATE_9216_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2187_l2190_l2197_DUPLICATE_ca71_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2187_l2190_l2197_DUPLICATE_ca71_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2187_l2190_l2197_DUPLICATE_ca71_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_2cd6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_2cd6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2187_l2174_l2197_DUPLICATE_e1af_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2187_l2174_l2197_DUPLICATE_e1af_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2187_l2174_l2197_DUPLICATE_e1af_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2174_c2_0f61_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2174_c2_0f61_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2174_c2_0f61_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2174_c2_0f61_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2197_c7_47bd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_e0af_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2197_c7_47bd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2174_c2_0f61] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2174_c2_0f61] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2174_c2_0f61] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2190_c7_8b8e] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond;
     t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output := t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2190_c7_8b8e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2174_c2_0f61] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2197_c7_47bd] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output := result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2197_c7_47bd] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_cond;
     t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output := t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2197_c7_47bd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2197_c7_47bd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_47bd_return_output;
     -- t16_high_MUX[uxn_opcodes_h_l2187_c7_85f5] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_cond;
     t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output := t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2190_c7_8b8e] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond;
     t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output := t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2190_c7_8b8e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2190_c7_8b8e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2190_c7_8b8e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2190_c7_8b8e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output := result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2187_c7_85f5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_8b8e_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2187_c7_85f5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output := result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2174_c2_0f61] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2174_c2_0f61] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_cond;
     t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output := t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2187_c7_85f5] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_cond;
     t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output := t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2187_c7_85f5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2187_c7_85f5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2187_c7_85f5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output;
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_85f5_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2174_c2_0f61] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2174_c2_0f61] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_cond;
     t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output := t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2174_c2_0f61] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2174_c2_0f61] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2174_c2_0f61] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output := result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output;

     -- Submodule level 5
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_ee25_uxn_opcodes_h_l2205_l2170_DUPLICATE_7b84 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ee25_uxn_opcodes_h_l2205_l2170_DUPLICATE_7b84_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_ee25(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_0f61_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ee25_uxn_opcodes_h_l2205_l2170_DUPLICATE_7b84_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ee25_uxn_opcodes_h_l2205_l2170_DUPLICATE_7b84_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
