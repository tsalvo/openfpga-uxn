-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 41
entity ldz_0CLK_a8170e34 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldz_0CLK_a8170e34;
architecture arch of ldz_0CLK_a8170e34 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1260_c6_31c9]
signal BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1260_c2_fd1b]
signal tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1260_c2_fd1b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1260_c2_fd1b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1260_c2_fd1b]
signal result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1260_c2_fd1b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1260_c2_fd1b]
signal result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1260_c2_fd1b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1260_c2_fd1b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1260_c2_fd1b]
signal t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1267_c11_60fe]
signal BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1267_c7_18eb]
signal tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1267_c7_18eb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1267_c7_18eb]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1267_c7_18eb]
signal result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1267_c7_18eb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1267_c7_18eb]
signal result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1267_c7_18eb]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1267_c7_18eb]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1267_c7_18eb]
signal t8_MUX_uxn_opcodes_h_l1267_c7_18eb_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1270_c30_96fc]
signal sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1272_c11_95f6]
signal BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1272_c7_a527]
signal tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1272_c7_a527]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1272_c7_a527]
signal result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1272_c7_a527]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1272_c7_a527]
signal result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1272_c7_a527]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1272_c7_a527]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1272_c7_a527]
signal t8_MUX_uxn_opcodes_h_l1272_c7_a527_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1272_c7_a527_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1278_c11_fa99]
signal BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1278_c7_f7cb]
signal tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1278_c7_f7cb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1278_c7_f7cb]
signal result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1278_c7_f7cb]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1278_c7_f7cb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1284_c11_0bd3]
signal BIN_OP_EQ_uxn_opcodes_h_l1284_c11_0bd3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1284_c11_0bd3_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1284_c11_0bd3_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1284_c7_5d92]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1284_c7_5d92]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_return_output : unsigned(0 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_44b7( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_stack_write := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9
BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_left,
BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_right,
BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b
tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond,
tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue,
tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse,
tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b
result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b
result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond,
result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b
result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b
result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b
result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output);

-- t8_MUX_uxn_opcodes_h_l1260_c2_fd1b
t8_MUX_uxn_opcodes_h_l1260_c2_fd1b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond,
t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue,
t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse,
t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe
BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_left,
BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_right,
BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb
tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_cond,
tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue,
tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse,
tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb
result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb
result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_cond,
result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb
result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb
result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_cond,
result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb
result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb
result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output);

-- t8_MUX_uxn_opcodes_h_l1267_c7_18eb
t8_MUX_uxn_opcodes_h_l1267_c7_18eb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1267_c7_18eb_cond,
t8_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue,
t8_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse,
t8_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc
sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_ins,
sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_x,
sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_y,
sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6
BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_left,
BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_right,
BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1272_c7_a527
tmp8_MUX_uxn_opcodes_h_l1272_c7_a527 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_cond,
tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue,
tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse,
tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527
result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527
result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_cond,
result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527
result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527
result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_cond,
result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527
result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_return_output);

-- t8_MUX_uxn_opcodes_h_l1272_c7_a527
t8_MUX_uxn_opcodes_h_l1272_c7_a527 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1272_c7_a527_cond,
t8_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue,
t8_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse,
t8_MUX_uxn_opcodes_h_l1272_c7_a527_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99
BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99_left,
BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99_right,
BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb
tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond,
tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue,
tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse,
tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb
result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb
result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond,
result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb
result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1284_c11_0bd3
BIN_OP_EQ_uxn_opcodes_h_l1284_c11_0bd3 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1284_c11_0bd3_left,
BIN_OP_EQ_uxn_opcodes_h_l1284_c11_0bd3_right,
BIN_OP_EQ_uxn_opcodes_h_l1284_c11_0bd3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92
result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92
result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_return_output,
 tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output,
 t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_return_output,
 tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output,
 t8_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output,
 sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_return_output,
 tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_return_output,
 t8_MUX_uxn_opcodes_h_l1272_c7_a527_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99_return_output,
 tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1284_c11_0bd3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1264_c3_8d97 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1268_c3_93e8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1272_c7_a527_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1267_c7_18eb_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1272_c7_a527_cond : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1275_c22_ec74_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1281_c3_a881 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c11_0bd3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c11_0bd3_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c11_0bd3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1272_l1260_DUPLICATE_9ef5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1272_l1267_l1260_DUPLICATE_8540_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1278_l1272_l1267_l1260_DUPLICATE_f288_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1267_l1260_DUPLICATE_f27a_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1284_l1272_l1267_l1260_DUPLICATE_7d0b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1284_l1278_l1272_l1267_DUPLICATE_546a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1278_l1272_DUPLICATE_4ab8_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_44b7_uxn_opcodes_h_l1289_l1256_DUPLICATE_214d_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c11_0bd3_right := to_unsigned(5, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1281_c3_a881 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1281_c3_a881;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1268_c3_93e8 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1268_c3_93e8;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1264_c3_8d97 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1264_c3_8d97;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c11_0bd3_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse := tmp8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1284_l1278_l1272_l1267_DUPLICATE_546a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1284_l1278_l1272_l1267_DUPLICATE_546a_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1278_c11_fa99] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99_left;
     BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99_return_output := BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1260_c6_31c9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_left;
     BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_return_output := BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1272_c11_95f6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_left;
     BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_return_output := BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_return_output;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1275_c22_ec74] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1275_c22_ec74_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1278_l1272_l1267_l1260_DUPLICATE_f288 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1278_l1272_l1267_l1260_DUPLICATE_f288_return_output := result.u8_value;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1278_l1272_DUPLICATE_4ab8 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1278_l1272_DUPLICATE_4ab8_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1267_c11_60fe] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_left;
     BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_return_output := BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1267_l1260_DUPLICATE_f27a LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1267_l1260_DUPLICATE_f27a_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1272_l1267_l1260_DUPLICATE_8540 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1272_l1267_l1260_DUPLICATE_8540_return_output := result.u16_value;

     -- sp_relative_shift[uxn_opcodes_h_l1270_c30_96fc] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_ins;
     sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_x;
     sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_return_output := sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1272_l1260_DUPLICATE_9ef5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1272_l1260_DUPLICATE_9ef5_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1284_l1272_l1267_l1260_DUPLICATE_7d0b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1284_l1272_l1267_l1260_DUPLICATE_7d0b_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1284_c11_0bd3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1284_c11_0bd3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c11_0bd3_left;
     BIN_OP_EQ_uxn_opcodes_h_l1284_c11_0bd3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c11_0bd3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c11_0bd3_return_output := BIN_OP_EQ_uxn_opcodes_h_l1284_c11_0bd3_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1260_c6_31c9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1267_c7_18eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1267_c11_60fe_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1272_c7_a527_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_95f6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_fa99_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c11_0bd3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1284_c11_0bd3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1275_c22_ec74_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1267_l1260_DUPLICATE_f27a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1267_l1260_DUPLICATE_f27a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1272_l1267_l1260_DUPLICATE_8540_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1272_l1267_l1260_DUPLICATE_8540_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1272_l1267_l1260_DUPLICATE_8540_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1284_l1278_l1272_l1267_DUPLICATE_546a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1284_l1278_l1272_l1267_DUPLICATE_546a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1284_l1278_l1272_l1267_DUPLICATE_546a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1284_l1278_l1272_l1267_DUPLICATE_546a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1272_l1260_DUPLICATE_9ef5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1272_l1260_DUPLICATE_9ef5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1284_l1272_l1267_l1260_DUPLICATE_7d0b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1284_l1272_l1267_l1260_DUPLICATE_7d0b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1284_l1272_l1267_l1260_DUPLICATE_7d0b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1284_l1272_l1267_l1260_DUPLICATE_7d0b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1278_l1272_DUPLICATE_4ab8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1278_l1272_DUPLICATE_4ab8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1278_l1272_l1267_l1260_DUPLICATE_f288_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1278_l1272_l1267_l1260_DUPLICATE_f288_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1278_l1272_l1267_l1260_DUPLICATE_f288_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1278_l1272_l1267_l1260_DUPLICATE_f288_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1270_c30_96fc_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1284_c7_5d92] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1284_c7_5d92] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1278_c7_f7cb] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output := result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1278_c7_f7cb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1278_c7_f7cb] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond;
     tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output := tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1267_c7_18eb] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output;

     -- t8_MUX[uxn_opcodes_h_l1272_c7_a527] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1272_c7_a527_cond <= VAR_t8_MUX_uxn_opcodes_h_l1272_c7_a527_cond;
     t8_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue;
     t8_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1272_c7_a527_return_output := t8_MUX_uxn_opcodes_h_l1272_c7_a527_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1272_c7_a527] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_return_output := result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1272_c7_a527] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1284_c7_5d92_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1272_c7_a527_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1284_c7_5d92_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1272_c7_a527_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1272_c7_a527_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1278_c7_f7cb] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1278_c7_f7cb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1272_c7_a527] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1260_c2_fd1b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1272_c7_a527] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_return_output := result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_return_output;

     -- t8_MUX[uxn_opcodes_h_l1267_c7_18eb] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1267_c7_18eb_cond <= VAR_t8_MUX_uxn_opcodes_h_l1267_c7_18eb_cond;
     t8_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue;
     t8_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output := t8_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1267_c7_18eb] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1267_c7_18eb] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output := result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1272_c7_a527] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_cond;
     tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_return_output := tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_f7cb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_a527_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_a527_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1272_c7_a527_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l1267_c7_18eb] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_cond;
     tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output := tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1267_c7_18eb] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output := result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1260_c2_fd1b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1272_c7_a527] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_return_output;

     -- t8_MUX[uxn_opcodes_h_l1260_c2_fd1b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond <= VAR_t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond;
     t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue;
     t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output := t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1272_c7_a527] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1260_c2_fd1b] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output := result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1267_c7_18eb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_a527_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_a527_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1267_c7_18eb] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1260_c2_fd1b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1260_c2_fd1b] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond;
     tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output := tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1260_c2_fd1b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1267_c7_18eb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1267_c7_18eb_return_output;
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1260_c2_fd1b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1260_c2_fd1b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_44b7_uxn_opcodes_h_l1289_l1256_DUPLICATE_214d LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_44b7_uxn_opcodes_h_l1289_l1256_DUPLICATE_214d_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_44b7(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1260_c2_fd1b_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_44b7_uxn_opcodes_h_l1289_l1256_DUPLICATE_214d_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_44b7_uxn_opcodes_h_l1289_l1256_DUPLICATE_214d_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
