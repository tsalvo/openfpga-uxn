-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 2
entity VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_0CLK_4b00ae23 is
port(
 ref_toks_0 : in uint8_t_80;
 var_dim_0 : in unsigned(6 downto 0);
 return_output : out unsigned(7 downto 0));
end VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_0CLK_4b00ae23;
architecture arch of VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_0CLK_4b00ae23 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- uint8_mux128[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2]
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_sel : unsigned(6 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in0 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in1 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in2 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in3 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in4 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in5 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in6 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in7 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in8 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in9 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in10 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in11 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in12 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in13 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in14 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in15 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in16 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in17 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in18 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in19 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in20 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in21 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in22 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in23 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in24 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in25 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in26 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in27 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in28 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in29 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in30 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in31 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in32 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in33 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in34 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in35 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in36 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in37 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in38 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in39 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in40 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in41 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in42 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in43 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in44 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in45 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in46 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in47 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in48 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in49 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in50 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in51 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in52 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in53 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in54 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in55 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in56 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in57 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in58 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in59 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in60 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in61 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in62 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in63 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in64 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in65 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in66 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in67 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in68 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in69 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in70 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in71 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in72 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in73 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in74 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in75 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in76 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in77 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in78 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in79 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in80 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in81 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in82 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in83 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in84 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in85 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in86 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in87 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in88 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in89 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in90 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in91 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in92 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in93 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in94 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in95 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in96 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in97 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in98 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in99 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in100 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in101 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in102 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in103 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in104 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in105 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in106 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in107 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in108 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in109 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in110 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in111 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in112 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in113 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in114 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in115 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in116 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in117 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in118 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in119 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in120 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in121 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in122 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in123 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in124 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in125 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in126 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in127 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_return_output : unsigned(7 downto 0);

function uint7_uint7_0( inp : unsigned;
 x : unsigned) return unsigned is

  --variable inp : unsigned(6 downto 0);
  --variable x : unsigned(6 downto 0);
  variable intermediate : unsigned(6 downto 0);
  variable return_output : unsigned(6 downto 0);

begin

    intermediate := (others => '0');
    intermediate(6 downto 0) := unsigned(inp);
    intermediate(6 downto 0) := x;
    
    return_output := intermediate(6 downto 0) ;
    
    return return_output;

end function;


begin

-- SUBMODULE INSTANCES 
-- uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2 : entity work.uint8_mux128_0CLK_9347d63d port map (
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_sel,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in0,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in1,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in2,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in3,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in4,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in5,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in6,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in7,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in8,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in9,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in10,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in11,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in12,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in13,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in14,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in15,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in16,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in17,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in18,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in19,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in20,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in21,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in22,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in23,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in24,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in25,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in26,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in27,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in28,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in29,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in30,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in31,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in32,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in33,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in34,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in35,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in36,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in37,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in38,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in39,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in40,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in41,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in42,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in43,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in44,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in45,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in46,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in47,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in48,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in49,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in50,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in51,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in52,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in53,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in54,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in55,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in56,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in57,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in58,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in59,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in60,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in61,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in62,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in63,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in64,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in65,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in66,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in67,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in68,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in69,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in70,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in71,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in72,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in73,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in74,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in75,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in76,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in77,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in78,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in79,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in80,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in81,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in82,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in83,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in84,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in85,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in86,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in87,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in88,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in89,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in90,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in91,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in92,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in93,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in94,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in95,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in96,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in97,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in98,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in99,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in100,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in101,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in102,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in103,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in104,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in105,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in106,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in107,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in108,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in109,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in110,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in111,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in112,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in113,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in114,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in115,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in116,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in117,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in118,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in119,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in120,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in121,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in122,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in123,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in124,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in125,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in126,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in127,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 ref_toks_0,
 var_dim_0,
 -- All submodule outputs
 uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_ref_toks_0 : uint8_t_80;
 variable VAR_var_dim_0 : unsigned(6 downto 0);
 variable VAR_return_output : unsigned(7 downto 0);
 variable VAR_base : uint8_t_80;
 variable VAR_ref_0 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_0_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l14_c10_c369_return_output : unsigned(7 downto 0);
 variable VAR_ref_1 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_1_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l16_c10_02db_return_output : unsigned(7 downto 0);
 variable VAR_ref_2 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_2_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l18_c10_a7d1_return_output : unsigned(7 downto 0);
 variable VAR_ref_3 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_3_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l20_c10_2ccf_return_output : unsigned(7 downto 0);
 variable VAR_ref_4 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_4_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l22_c10_19e4_return_output : unsigned(7 downto 0);
 variable VAR_ref_5 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_5_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l24_c10_0618_return_output : unsigned(7 downto 0);
 variable VAR_ref_6 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_6_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l26_c10_357e_return_output : unsigned(7 downto 0);
 variable VAR_ref_7 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_7_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l28_c10_348f_return_output : unsigned(7 downto 0);
 variable VAR_ref_8 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_8_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l30_c10_8a3b_return_output : unsigned(7 downto 0);
 variable VAR_ref_9 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_9_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l32_c10_be34_return_output : unsigned(7 downto 0);
 variable VAR_ref_10 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_10_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l34_c11_6fc1_return_output : unsigned(7 downto 0);
 variable VAR_ref_11 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_11_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l36_c11_ad43_return_output : unsigned(7 downto 0);
 variable VAR_ref_12 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_12_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l38_c11_ccb7_return_output : unsigned(7 downto 0);
 variable VAR_ref_13 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_13_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l40_c11_d2d2_return_output : unsigned(7 downto 0);
 variable VAR_ref_14 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_14_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l42_c11_89b8_return_output : unsigned(7 downto 0);
 variable VAR_ref_15 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_15_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l44_c11_be8b_return_output : unsigned(7 downto 0);
 variable VAR_ref_16 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_16_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l46_c11_14bf_return_output : unsigned(7 downto 0);
 variable VAR_ref_17 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_17_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l48_c11_c516_return_output : unsigned(7 downto 0);
 variable VAR_ref_18 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_18_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l50_c11_d116_return_output : unsigned(7 downto 0);
 variable VAR_ref_19 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_19_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l52_c11_2334_return_output : unsigned(7 downto 0);
 variable VAR_ref_20 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_20_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l54_c11_a600_return_output : unsigned(7 downto 0);
 variable VAR_ref_21 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_21_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l56_c11_09c6_return_output : unsigned(7 downto 0);
 variable VAR_ref_22 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_22_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l58_c11_a4bb_return_output : unsigned(7 downto 0);
 variable VAR_ref_23 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_23_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l60_c11_fe80_return_output : unsigned(7 downto 0);
 variable VAR_ref_24 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_24_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l62_c11_5300_return_output : unsigned(7 downto 0);
 variable VAR_ref_25 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_25_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l64_c11_8cbd_return_output : unsigned(7 downto 0);
 variable VAR_ref_26 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_26_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l66_c11_749a_return_output : unsigned(7 downto 0);
 variable VAR_ref_27 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_27_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l68_c11_bd2e_return_output : unsigned(7 downto 0);
 variable VAR_ref_28 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_28_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l70_c11_14ca_return_output : unsigned(7 downto 0);
 variable VAR_ref_29 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_29_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l72_c11_438c_return_output : unsigned(7 downto 0);
 variable VAR_ref_30 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_30_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l74_c11_e26a_return_output : unsigned(7 downto 0);
 variable VAR_ref_31 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_31_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l76_c11_2bbd_return_output : unsigned(7 downto 0);
 variable VAR_ref_32 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_32_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l78_c11_3450_return_output : unsigned(7 downto 0);
 variable VAR_ref_33 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_33_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l80_c11_da79_return_output : unsigned(7 downto 0);
 variable VAR_ref_34 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_34_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l82_c11_de59_return_output : unsigned(7 downto 0);
 variable VAR_ref_35 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_35_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l84_c11_83cd_return_output : unsigned(7 downto 0);
 variable VAR_ref_36 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_36_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l86_c11_5632_return_output : unsigned(7 downto 0);
 variable VAR_ref_37 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_37_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l88_c11_34a2_return_output : unsigned(7 downto 0);
 variable VAR_ref_38 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_38_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l90_c11_7b08_return_output : unsigned(7 downto 0);
 variable VAR_ref_39 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_39_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l92_c11_5674_return_output : unsigned(7 downto 0);
 variable VAR_ref_40 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_40_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l94_c11_17f2_return_output : unsigned(7 downto 0);
 variable VAR_ref_41 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_41_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l96_c11_e556_return_output : unsigned(7 downto 0);
 variable VAR_ref_42 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_42_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l98_c11_067a_return_output : unsigned(7 downto 0);
 variable VAR_ref_43 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_43_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l100_c11_c543_return_output : unsigned(7 downto 0);
 variable VAR_ref_44 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_44_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l102_c11_dc88_return_output : unsigned(7 downto 0);
 variable VAR_ref_45 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_45_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l104_c11_5ee7_return_output : unsigned(7 downto 0);
 variable VAR_ref_46 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_46_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l106_c11_7288_return_output : unsigned(7 downto 0);
 variable VAR_ref_47 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_47_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l108_c11_fb1f_return_output : unsigned(7 downto 0);
 variable VAR_ref_48 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_48_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l110_c11_89c3_return_output : unsigned(7 downto 0);
 variable VAR_ref_49 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_49_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l112_c11_ae5c_return_output : unsigned(7 downto 0);
 variable VAR_ref_50 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_50_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l114_c11_25eb_return_output : unsigned(7 downto 0);
 variable VAR_ref_51 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_51_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l116_c11_49c5_return_output : unsigned(7 downto 0);
 variable VAR_ref_52 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_52_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l118_c11_4de9_return_output : unsigned(7 downto 0);
 variable VAR_ref_53 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_53_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l120_c11_0207_return_output : unsigned(7 downto 0);
 variable VAR_ref_54 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_54_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l122_c11_4729_return_output : unsigned(7 downto 0);
 variable VAR_ref_55 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_55_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l124_c11_92df_return_output : unsigned(7 downto 0);
 variable VAR_ref_56 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_56_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l126_c11_e0b6_return_output : unsigned(7 downto 0);
 variable VAR_ref_57 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_57_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l128_c11_628c_return_output : unsigned(7 downto 0);
 variable VAR_ref_58 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_58_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l130_c11_31ac_return_output : unsigned(7 downto 0);
 variable VAR_ref_59 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_59_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l132_c11_4a25_return_output : unsigned(7 downto 0);
 variable VAR_ref_60 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_60_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l134_c11_20a3_return_output : unsigned(7 downto 0);
 variable VAR_ref_61 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_61_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l136_c11_3776_return_output : unsigned(7 downto 0);
 variable VAR_ref_62 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_62_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l138_c11_6592_return_output : unsigned(7 downto 0);
 variable VAR_ref_63 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_63_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l140_c11_fe1a_return_output : unsigned(7 downto 0);
 variable VAR_ref_64 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_64_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l142_c11_d869_return_output : unsigned(7 downto 0);
 variable VAR_ref_65 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_65_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l144_c11_f34d_return_output : unsigned(7 downto 0);
 variable VAR_ref_66 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_66_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l146_c11_5734_return_output : unsigned(7 downto 0);
 variable VAR_ref_67 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_67_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l148_c11_5797_return_output : unsigned(7 downto 0);
 variable VAR_ref_68 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_68_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l150_c11_38e6_return_output : unsigned(7 downto 0);
 variable VAR_ref_69 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_69_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l152_c11_9f83_return_output : unsigned(7 downto 0);
 variable VAR_ref_70 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_70_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l154_c11_d8d3_return_output : unsigned(7 downto 0);
 variable VAR_ref_71 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_71_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l156_c11_0e0a_return_output : unsigned(7 downto 0);
 variable VAR_ref_72 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_72_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l158_c11_8a55_return_output : unsigned(7 downto 0);
 variable VAR_ref_73 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_73_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l160_c11_a527_return_output : unsigned(7 downto 0);
 variable VAR_ref_74 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_74_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l162_c11_ea69_return_output : unsigned(7 downto 0);
 variable VAR_ref_75 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_75_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l164_c11_686b_return_output : unsigned(7 downto 0);
 variable VAR_ref_76 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_76_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l166_c11_c767_return_output : unsigned(7 downto 0);
 variable VAR_ref_77 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_77_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l168_c11_d44f_return_output : unsigned(7 downto 0);
 variable VAR_ref_78 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_78_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l170_c11_3b86_return_output : unsigned(7 downto 0);
 variable VAR_ref_79 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output : unsigned(7 downto 0);
 variable VAR_sel : unsigned(6 downto 0);
 variable VAR_sel_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l175_c2_0829 : unsigned(6 downto 0);
 variable VAR_uint7_uint7_0_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l176_c8_153f_return_output : unsigned(6 downto 0);
 variable VAR_rv : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_sel : unsigned(6 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in0 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in1 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in2 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in3 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in4 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in5 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in6 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in7 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in8 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in9 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in10 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in11 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in12 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in13 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in14 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in15 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in16 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in17 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in18 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in19 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in20 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in21 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in22 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in23 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in24 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in25 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in26 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in27 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in28 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in29 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in30 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in31 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in32 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in33 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in34 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in35 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in36 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in37 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in38 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in39 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in40 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in41 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in42 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in43 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in44 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in45 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in46 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in47 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in48 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in49 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in50 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in51 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in52 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in53 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in54 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in55 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in56 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in57 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in58 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in59 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in60 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in61 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in62 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in63 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in64 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in65 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in66 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in67 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in68 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in69 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in70 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in71 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in72 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in73 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in74 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in75 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in76 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in77 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in78 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in79 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in80 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in81 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in82 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in83 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in84 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in85 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in86 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in87 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in88 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in89 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in90 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in91 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in92 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in93 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in94 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in95 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in96 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in97 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in98 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in99 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in100 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in101 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in102 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in103 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in104 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in105 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in106 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in107 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in108 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in109 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in110 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in111 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in112 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in113 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in114 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in115 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in116 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in117 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in118 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in119 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in120 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in121 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in122 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in123 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in124 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in125 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in126 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in127 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_return_output : unsigned(7 downto 0);
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sel_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l175_c2_0829 := resize(to_unsigned(0, 1), 7);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_ref_toks_0 := ref_toks_0;
     VAR_var_dim_0 := var_dim_0;

     -- Submodule level 0
     -- CONST_REF_RD_uint8_t_uint8_t_80_37_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l88_c11_34a2] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_37_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l88_c11_34a2_return_output := VAR_ref_toks_0(37);

     -- CONST_REF_RD_uint8_t_uint8_t_80_74_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l162_c11_ea69] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_74_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l162_c11_ea69_return_output := VAR_ref_toks_0(74);

     -- CONST_REF_RD_uint8_t_uint8_t_80_9_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l32_c10_be34] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_9_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l32_c10_be34_return_output := VAR_ref_toks_0(9);

     -- CONST_REF_RD_uint8_t_uint8_t_80_64_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l142_c11_d869] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_64_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l142_c11_d869_return_output := VAR_ref_toks_0(64);

     -- CONST_REF_RD_uint8_t_uint8_t_80_17_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l48_c11_c516] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_17_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l48_c11_c516_return_output := VAR_ref_toks_0(17);

     -- CONST_REF_RD_uint8_t_uint8_t_80_65_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l144_c11_f34d] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_65_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l144_c11_f34d_return_output := VAR_ref_toks_0(65);

     -- CONST_REF_RD_uint8_t_uint8_t_80_72_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l158_c11_8a55] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_72_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l158_c11_8a55_return_output := VAR_ref_toks_0(72);

     -- CONST_REF_RD_uint8_t_uint8_t_80_12_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l38_c11_ccb7] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_12_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l38_c11_ccb7_return_output := VAR_ref_toks_0(12);

     -- CONST_REF_RD_uint8_t_uint8_t_80_56_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l126_c11_e0b6] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_56_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l126_c11_e0b6_return_output := VAR_ref_toks_0(56);

     -- CONST_REF_RD_uint8_t_uint8_t_80_69_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l152_c11_9f83] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_69_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l152_c11_9f83_return_output := VAR_ref_toks_0(69);

     -- CONST_REF_RD_uint8_t_uint8_t_80_24_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l62_c11_5300] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_24_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l62_c11_5300_return_output := VAR_ref_toks_0(24);

     -- CONST_REF_RD_uint8_t_uint8_t_80_26_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l66_c11_749a] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_26_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l66_c11_749a_return_output := VAR_ref_toks_0(26);

     -- CONST_REF_RD_uint8_t_uint8_t_80_79_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output := VAR_ref_toks_0(79);

     -- CONST_REF_RD_uint8_t_uint8_t_80_60_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l134_c11_20a3] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_60_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l134_c11_20a3_return_output := VAR_ref_toks_0(60);

     -- CONST_REF_RD_uint8_t_uint8_t_80_33_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l80_c11_da79] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_33_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l80_c11_da79_return_output := VAR_ref_toks_0(33);

     -- CONST_REF_RD_uint8_t_uint8_t_80_13_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l40_c11_d2d2] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_13_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l40_c11_d2d2_return_output := VAR_ref_toks_0(13);

     -- CONST_REF_RD_uint8_t_uint8_t_80_71_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l156_c11_0e0a] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_71_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l156_c11_0e0a_return_output := VAR_ref_toks_0(71);

     -- CONST_REF_RD_uint8_t_uint8_t_80_42_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l98_c11_067a] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_42_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l98_c11_067a_return_output := VAR_ref_toks_0(42);

     -- CONST_REF_RD_uint8_t_uint8_t_80_55_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l124_c11_92df] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_55_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l124_c11_92df_return_output := VAR_ref_toks_0(55);

     -- CONST_REF_RD_uint8_t_uint8_t_80_43_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l100_c11_c543] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_43_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l100_c11_c543_return_output := VAR_ref_toks_0(43);

     -- CONST_REF_RD_uint8_t_uint8_t_80_15_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l44_c11_be8b] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_15_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l44_c11_be8b_return_output := VAR_ref_toks_0(15);

     -- CONST_REF_RD_uint8_t_uint8_t_80_27_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l68_c11_bd2e] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_27_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l68_c11_bd2e_return_output := VAR_ref_toks_0(27);

     -- CONST_REF_RD_uint8_t_uint8_t_80_59_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l132_c11_4a25] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_59_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l132_c11_4a25_return_output := VAR_ref_toks_0(59);

     -- CONST_REF_RD_uint8_t_uint8_t_80_16_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l46_c11_14bf] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_16_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l46_c11_14bf_return_output := VAR_ref_toks_0(16);

     -- CONST_REF_RD_uint8_t_uint8_t_80_22_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l58_c11_a4bb] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_22_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l58_c11_a4bb_return_output := VAR_ref_toks_0(22);

     -- CONST_REF_RD_uint8_t_uint8_t_80_36_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l86_c11_5632] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_36_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l86_c11_5632_return_output := VAR_ref_toks_0(36);

     -- CONST_REF_RD_uint8_t_uint8_t_80_0_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l14_c10_c369] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_0_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l14_c10_c369_return_output := VAR_ref_toks_0(0);

     -- CONST_REF_RD_uint8_t_uint8_t_80_20_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l54_c11_a600] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_20_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l54_c11_a600_return_output := VAR_ref_toks_0(20);

     -- CONST_REF_RD_uint8_t_uint8_t_80_29_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l72_c11_438c] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_29_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l72_c11_438c_return_output := VAR_ref_toks_0(29);

     -- CONST_REF_RD_uint8_t_uint8_t_80_57_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l128_c11_628c] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_57_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l128_c11_628c_return_output := VAR_ref_toks_0(57);

     -- CONST_REF_RD_uint8_t_uint8_t_80_61_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l136_c11_3776] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_61_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l136_c11_3776_return_output := VAR_ref_toks_0(61);

     -- CONST_REF_RD_uint8_t_uint8_t_80_53_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l120_c11_0207] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_53_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l120_c11_0207_return_output := VAR_ref_toks_0(53);

     -- CONST_REF_RD_uint8_t_uint8_t_80_52_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l118_c11_4de9] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_52_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l118_c11_4de9_return_output := VAR_ref_toks_0(52);

     -- CONST_REF_RD_uint8_t_uint8_t_80_70_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l154_c11_d8d3] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_70_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l154_c11_d8d3_return_output := VAR_ref_toks_0(70);

     -- CONST_REF_RD_uint8_t_uint8_t_80_32_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l78_c11_3450] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_32_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l78_c11_3450_return_output := VAR_ref_toks_0(32);

     -- CONST_REF_RD_uint8_t_uint8_t_80_51_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l116_c11_49c5] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_51_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l116_c11_49c5_return_output := VAR_ref_toks_0(51);

     -- CONST_REF_RD_uint8_t_uint8_t_80_21_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l56_c11_09c6] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_21_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l56_c11_09c6_return_output := VAR_ref_toks_0(21);

     -- CONST_REF_RD_uint8_t_uint8_t_80_28_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l70_c11_14ca] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_28_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l70_c11_14ca_return_output := VAR_ref_toks_0(28);

     -- uint7_uint7_0[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l176_c8_153f] LATENCY=0
     VAR_uint7_uint7_0_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l176_c8_153f_return_output := uint7_uint7_0(
     VAR_sel_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l175_c2_0829,
     VAR_var_dim_0);

     -- CONST_REF_RD_uint8_t_uint8_t_80_5_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l24_c10_0618] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_5_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l24_c10_0618_return_output := VAR_ref_toks_0(5);

     -- CONST_REF_RD_uint8_t_uint8_t_80_39_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l92_c11_5674] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_39_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l92_c11_5674_return_output := VAR_ref_toks_0(39);

     -- CONST_REF_RD_uint8_t_uint8_t_80_1_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l16_c10_02db] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_1_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l16_c10_02db_return_output := VAR_ref_toks_0(1);

     -- CONST_REF_RD_uint8_t_uint8_t_80_38_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l90_c11_7b08] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_38_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l90_c11_7b08_return_output := VAR_ref_toks_0(38);

     -- CONST_REF_RD_uint8_t_uint8_t_80_10_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l34_c11_6fc1] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_10_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l34_c11_6fc1_return_output := VAR_ref_toks_0(10);

     -- CONST_REF_RD_uint8_t_uint8_t_80_3_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l20_c10_2ccf] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_3_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l20_c10_2ccf_return_output := VAR_ref_toks_0(3);

     -- CONST_REF_RD_uint8_t_uint8_t_80_25_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l64_c11_8cbd] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_25_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l64_c11_8cbd_return_output := VAR_ref_toks_0(25);

     -- CONST_REF_RD_uint8_t_uint8_t_80_18_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l50_c11_d116] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_18_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l50_c11_d116_return_output := VAR_ref_toks_0(18);

     -- CONST_REF_RD_uint8_t_uint8_t_80_77_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l168_c11_d44f] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_77_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l168_c11_d44f_return_output := VAR_ref_toks_0(77);

     -- CONST_REF_RD_uint8_t_uint8_t_80_62_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l138_c11_6592] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_62_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l138_c11_6592_return_output := VAR_ref_toks_0(62);

     -- CONST_REF_RD_uint8_t_uint8_t_80_49_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l112_c11_ae5c] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_49_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l112_c11_ae5c_return_output := VAR_ref_toks_0(49);

     -- CONST_REF_RD_uint8_t_uint8_t_80_46_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l106_c11_7288] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_46_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l106_c11_7288_return_output := VAR_ref_toks_0(46);

     -- CONST_REF_RD_uint8_t_uint8_t_80_14_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l42_c11_89b8] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_14_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l42_c11_89b8_return_output := VAR_ref_toks_0(14);

     -- CONST_REF_RD_uint8_t_uint8_t_80_31_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l76_c11_2bbd] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_31_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l76_c11_2bbd_return_output := VAR_ref_toks_0(31);

     -- CONST_REF_RD_uint8_t_uint8_t_80_47_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l108_c11_fb1f] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_47_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l108_c11_fb1f_return_output := VAR_ref_toks_0(47);

     -- CONST_REF_RD_uint8_t_uint8_t_80_34_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l82_c11_de59] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_34_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l82_c11_de59_return_output := VAR_ref_toks_0(34);

     -- CONST_REF_RD_uint8_t_uint8_t_80_67_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l148_c11_5797] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_67_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l148_c11_5797_return_output := VAR_ref_toks_0(67);

     -- CONST_REF_RD_uint8_t_uint8_t_80_66_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l146_c11_5734] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_66_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l146_c11_5734_return_output := VAR_ref_toks_0(66);

     -- CONST_REF_RD_uint8_t_uint8_t_80_78_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l170_c11_3b86] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_78_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l170_c11_3b86_return_output := VAR_ref_toks_0(78);

     -- CONST_REF_RD_uint8_t_uint8_t_80_2_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l18_c10_a7d1] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_2_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l18_c10_a7d1_return_output := VAR_ref_toks_0(2);

     -- CONST_REF_RD_uint8_t_uint8_t_80_54_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l122_c11_4729] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_54_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l122_c11_4729_return_output := VAR_ref_toks_0(54);

     -- CONST_REF_RD_uint8_t_uint8_t_80_23_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l60_c11_fe80] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_23_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l60_c11_fe80_return_output := VAR_ref_toks_0(23);

     -- CONST_REF_RD_uint8_t_uint8_t_80_58_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l130_c11_31ac] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_58_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l130_c11_31ac_return_output := VAR_ref_toks_0(58);

     -- CONST_REF_RD_uint8_t_uint8_t_80_30_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l74_c11_e26a] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_30_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l74_c11_e26a_return_output := VAR_ref_toks_0(30);

     -- CONST_REF_RD_uint8_t_uint8_t_80_7_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l28_c10_348f] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_7_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l28_c10_348f_return_output := VAR_ref_toks_0(7);

     -- CONST_REF_RD_uint8_t_uint8_t_80_48_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l110_c11_89c3] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_48_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l110_c11_89c3_return_output := VAR_ref_toks_0(48);

     -- CONST_REF_RD_uint8_t_uint8_t_80_73_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l160_c11_a527] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_73_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l160_c11_a527_return_output := VAR_ref_toks_0(73);

     -- CONST_REF_RD_uint8_t_uint8_t_80_8_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l30_c10_8a3b] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_8_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l30_c10_8a3b_return_output := VAR_ref_toks_0(8);

     -- CONST_REF_RD_uint8_t_uint8_t_80_45_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l104_c11_5ee7] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_45_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l104_c11_5ee7_return_output := VAR_ref_toks_0(45);

     -- CONST_REF_RD_uint8_t_uint8_t_80_63_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l140_c11_fe1a] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_63_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l140_c11_fe1a_return_output := VAR_ref_toks_0(63);

     -- CONST_REF_RD_uint8_t_uint8_t_80_50_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l114_c11_25eb] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_50_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l114_c11_25eb_return_output := VAR_ref_toks_0(50);

     -- CONST_REF_RD_uint8_t_uint8_t_80_75_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l164_c11_686b] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_75_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l164_c11_686b_return_output := VAR_ref_toks_0(75);

     -- CONST_REF_RD_uint8_t_uint8_t_80_44_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l102_c11_dc88] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_44_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l102_c11_dc88_return_output := VAR_ref_toks_0(44);

     -- CONST_REF_RD_uint8_t_uint8_t_80_68_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l150_c11_38e6] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_68_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l150_c11_38e6_return_output := VAR_ref_toks_0(68);

     -- CONST_REF_RD_uint8_t_uint8_t_80_76_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l166_c11_c767] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_76_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l166_c11_c767_return_output := VAR_ref_toks_0(76);

     -- CONST_REF_RD_uint8_t_uint8_t_80_19_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l52_c11_2334] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_19_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l52_c11_2334_return_output := VAR_ref_toks_0(19);

     -- CONST_REF_RD_uint8_t_uint8_t_80_6_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l26_c10_357e] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_6_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l26_c10_357e_return_output := VAR_ref_toks_0(6);

     -- CONST_REF_RD_uint8_t_uint8_t_80_35_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l84_c11_83cd] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_35_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l84_c11_83cd_return_output := VAR_ref_toks_0(35);

     -- CONST_REF_RD_uint8_t_uint8_t_80_40_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l94_c11_17f2] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_40_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l94_c11_17f2_return_output := VAR_ref_toks_0(40);

     -- CONST_REF_RD_uint8_t_uint8_t_80_41_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l96_c11_e556] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_41_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l96_c11_e556_return_output := VAR_ref_toks_0(41);

     -- CONST_REF_RD_uint8_t_uint8_t_80_11_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l36_c11_ad43] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_11_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l36_c11_ad43_return_output := VAR_ref_toks_0(11);

     -- CONST_REF_RD_uint8_t_uint8_t_80_4_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l22_c10_19e4] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_4_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l22_c10_19e4_return_output := VAR_ref_toks_0(4);

     -- Submodule level 1
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in0 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_0_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l14_c10_c369_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in10 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_10_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l34_c11_6fc1_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in11 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_11_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l36_c11_ad43_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in12 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_12_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l38_c11_ccb7_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in13 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_13_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l40_c11_d2d2_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in14 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_14_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l42_c11_89b8_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in15 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_15_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l44_c11_be8b_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in16 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_16_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l46_c11_14bf_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in17 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_17_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l48_c11_c516_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in18 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_18_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l50_c11_d116_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in19 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_19_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l52_c11_2334_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in1 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_1_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l16_c10_02db_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in20 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_20_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l54_c11_a600_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in21 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_21_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l56_c11_09c6_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in22 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_22_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l58_c11_a4bb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in23 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_23_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l60_c11_fe80_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in24 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_24_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l62_c11_5300_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in25 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_25_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l64_c11_8cbd_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in26 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_26_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l66_c11_749a_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in27 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_27_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l68_c11_bd2e_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in28 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_28_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l70_c11_14ca_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in29 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_29_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l72_c11_438c_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in2 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_2_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l18_c10_a7d1_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in30 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_30_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l74_c11_e26a_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in31 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_31_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l76_c11_2bbd_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in32 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_32_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l78_c11_3450_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in33 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_33_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l80_c11_da79_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in34 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_34_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l82_c11_de59_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in35 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_35_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l84_c11_83cd_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in36 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_36_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l86_c11_5632_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in37 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_37_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l88_c11_34a2_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in38 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_38_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l90_c11_7b08_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in39 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_39_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l92_c11_5674_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in3 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_3_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l20_c10_2ccf_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in40 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_40_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l94_c11_17f2_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in41 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_41_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l96_c11_e556_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in42 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_42_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l98_c11_067a_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in43 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_43_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l100_c11_c543_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in44 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_44_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l102_c11_dc88_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in45 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_45_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l104_c11_5ee7_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in46 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_46_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l106_c11_7288_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in47 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_47_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l108_c11_fb1f_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in48 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_48_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l110_c11_89c3_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in49 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_49_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l112_c11_ae5c_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in4 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_4_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l22_c10_19e4_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in50 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_50_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l114_c11_25eb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in51 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_51_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l116_c11_49c5_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in52 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_52_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l118_c11_4de9_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in53 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_53_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l120_c11_0207_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in54 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_54_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l122_c11_4729_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in55 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_55_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l124_c11_92df_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in56 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_56_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l126_c11_e0b6_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in57 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_57_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l128_c11_628c_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in58 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_58_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l130_c11_31ac_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in59 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_59_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l132_c11_4a25_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in5 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_5_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l24_c10_0618_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in60 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_60_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l134_c11_20a3_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in61 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_61_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l136_c11_3776_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in62 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_62_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l138_c11_6592_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in63 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_63_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l140_c11_fe1a_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in64 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_64_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l142_c11_d869_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in65 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_65_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l144_c11_f34d_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in66 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_66_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l146_c11_5734_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in67 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_67_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l148_c11_5797_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in68 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_68_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l150_c11_38e6_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in69 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_69_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l152_c11_9f83_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in6 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_6_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l26_c10_357e_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in70 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_70_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l154_c11_d8d3_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in71 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_71_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l156_c11_0e0a_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in72 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_72_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l158_c11_8a55_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in73 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_73_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l160_c11_a527_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in74 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_74_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l162_c11_ea69_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in75 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_75_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l164_c11_686b_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in76 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_76_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l166_c11_c767_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in77 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_77_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l168_c11_d44f_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in78 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_78_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l170_c11_3b86_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in100 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in101 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in102 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in103 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in104 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in105 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in106 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in107 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in108 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in109 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in110 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in111 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in112 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in113 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in114 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in115 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in116 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in117 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in118 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in119 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in120 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in121 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in122 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in123 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in124 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in125 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in126 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in127 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in79 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in80 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in81 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in82 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in83 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in84 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in85 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in86 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in87 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in88 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in89 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in90 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in91 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in92 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in93 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in94 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in95 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in96 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in97 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in98 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in99 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_ec09_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in7 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_7_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l28_c10_348f_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in8 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_8_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l30_c10_8a3b_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in9 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_9_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l32_c10_be34_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_sel := VAR_uint7_uint7_0_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l176_c8_153f_return_output;
     -- uint8_mux128[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2] LATENCY=0
     -- Inputs
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_sel <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_sel;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in0 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in0;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in1 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in1;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in2 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in2;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in3 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in3;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in4 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in4;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in5 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in5;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in6 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in6;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in7 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in7;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in8 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in8;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in9 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in9;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in10 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in10;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in11 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in11;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in12 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in12;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in13 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in13;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in14 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in14;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in15 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in15;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in16 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in16;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in17 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in17;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in18 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in18;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in19 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in19;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in20 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in20;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in21 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in21;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in22 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in22;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in23 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in23;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in24 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in24;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in25 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in25;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in26 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in26;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in27 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in27;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in28 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in28;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in29 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in29;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in30 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in30;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in31 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in31;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in32 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in32;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in33 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in33;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in34 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in34;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in35 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in35;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in36 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in36;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in37 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in37;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in38 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in38;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in39 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in39;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in40 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in40;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in41 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in41;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in42 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in42;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in43 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in43;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in44 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in44;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in45 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in45;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in46 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in46;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in47 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in47;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in48 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in48;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in49 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in49;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in50 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in50;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in51 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in51;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in52 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in52;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in53 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in53;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in54 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in54;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in55 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in55;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in56 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in56;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in57 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in57;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in58 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in58;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in59 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in59;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in60 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in60;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in61 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in61;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in62 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in62;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in63 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in63;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in64 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in64;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in65 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in65;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in66 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in66;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in67 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in67;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in68 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in68;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in69 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in69;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in70 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in70;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in71 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in71;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in72 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in72;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in73 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in73;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in74 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in74;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in75 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in75;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in76 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in76;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in77 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in77;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in78 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in78;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in79 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in79;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in80 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in80;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in81 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in81;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in82 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in82;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in83 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in83;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in84 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in84;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in85 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in85;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in86 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in86;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in87 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in87;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in88 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in88;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in89 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in89;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in90 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in90;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in91 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in91;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in92 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in92;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in93 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in93;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in94 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in94;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in95 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in95;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in96 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in96;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in97 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in97;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in98 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in98;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in99 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in99;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in100 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in100;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in101 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in101;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in102 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in102;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in103 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in103;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in104 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in104;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in105 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in105;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in106 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in106;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in107 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in107;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in108 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in108;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in109 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in109;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in110 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in110;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in111 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in111;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in112 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in112;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in113 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in113;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in114 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in114;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in115 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in115;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in116 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in116;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in117 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in117;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in118 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in118;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in119 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in119;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in120 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in120;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in121 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in121;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in122 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in122;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in123 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in123;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in124 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in124;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in125 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in125;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in126 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in126;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in127 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_in127;
     -- Outputs
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_return_output := uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_return_output;

     -- Submodule level 2
     VAR_return_output := VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_10e2_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
