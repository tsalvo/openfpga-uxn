-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity sth2_0CLK_55b6500a is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sth2_0CLK_55b6500a;
architecture arch of sth2_0CLK_55b6500a is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2420_c6_fee1]
signal BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2420_c2_fc3f]
signal t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2420_c2_fc3f]
signal t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2420_c2_fc3f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2420_c2_fc3f]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2420_c2_fc3f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2420_c2_fc3f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2420_c2_fc3f]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2420_c2_fc3f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2420_c2_fc3f]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2420_c2_fc3f]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2420_c2_fc3f]
signal result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2433_c11_1b72]
signal BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2433_c7_fcec]
signal t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2433_c7_fcec]
signal t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2433_c7_fcec]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2433_c7_fcec]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2433_c7_fcec]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2433_c7_fcec]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2433_c7_fcec]
signal result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2433_c7_fcec]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2436_c11_299c]
signal BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2436_c7_07dd]
signal t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2436_c7_07dd]
signal t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2436_c7_07dd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2436_c7_07dd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2436_c7_07dd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2436_c7_07dd]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2436_c7_07dd]
signal result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2436_c7_07dd]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2438_c30_3f27]
signal sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2440_c11_ea1d]
signal BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2440_c7_fedf]
signal t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2440_c7_fedf]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2440_c7_fedf]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2440_c7_fedf]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2440_c7_fedf]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2440_c7_fedf]
signal result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2440_c7_fedf]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2448_c11_184a]
signal BIN_OP_EQ_uxn_opcodes_h_l2448_c11_184a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2448_c11_184a_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2448_c11_184a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2448_c7_decb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2448_c7_decb]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2448_c7_decb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2448_c7_decb]
signal result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_04b4( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.is_stack_index_flipped := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.u8_value := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1
BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_left,
BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_right,
BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f
t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond,
t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue,
t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse,
t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f
t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond,
t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue,
t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse,
t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f
result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f
result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f
result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f
result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f
result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f
result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72
BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_left,
BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_right,
BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec
t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_cond,
t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue,
t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse,
t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec
t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_cond,
t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue,
t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse,
t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec
result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec
result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec
result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec
result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_cond,
result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c
BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_left,
BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_right,
BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd
t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_cond,
t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue,
t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse,
t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd
t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_cond,
t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue,
t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse,
t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd
result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd
result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd
result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd
result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_cond,
result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27
sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_ins,
sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_x,
sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_y,
sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d
BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_left,
BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_right,
BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf
t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_cond,
t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue,
t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse,
t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf
result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf
result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf
result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf
result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_cond,
result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2448_c11_184a
BIN_OP_EQ_uxn_opcodes_h_l2448_c11_184a : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2448_c11_184a_left,
BIN_OP_EQ_uxn_opcodes_h_l2448_c11_184a_right,
BIN_OP_EQ_uxn_opcodes_h_l2448_c11_184a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb
result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb
result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb
result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_cond,
result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_return_output,
 t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output,
 t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_return_output,
 t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output,
 t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_return_output,
 t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output,
 t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output,
 sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_return_output,
 t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2448_c11_184a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2420_c2_fc3f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2430_c3_bb63 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2425_c3_0f2c : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2420_c2_fc3f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2420_c2_fc3f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2434_c3_58d1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2443_c3_53c9 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2445_c3_536a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c11_184a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c11_184a_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c11_184a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2449_c3_8719 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2450_c3_c149 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2420_l2433_l2448_l2436_DUPLICATE_a81a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2433_l2448_DUPLICATE_4c62_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2440_l2433_l2448_l2436_DUPLICATE_87de_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2440_l2433_l2436_DUPLICATE_7f8b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2440_l2433_l2436_DUPLICATE_27db_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2448_l2436_DUPLICATE_28e9_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2455_l2416_DUPLICATE_84a1_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c11_184a_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2445_c3_536a := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2445_c3_536a;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_right := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2449_c3_8719 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2449_c3_8719;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2443_c3_53c9 := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2443_c3_53c9;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_y := resize(to_signed(-2, 3), 4);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2434_c3_58d1 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2434_c3_58d1;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2450_c3_c149 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2450_c3_c149;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2425_c3_0f2c := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2425_c3_0f2c;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2430_c3_bb63 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2430_c3_bb63;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_right := to_unsigned(2, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c11_184a_left := VAR_phase;
     VAR_t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue := VAR_previous_stack_read;
     VAR_t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse := t16_high;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse := t16_low;
     -- BIN_OP_EQ[uxn_opcodes_h_l2440_c11_ea1d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_left;
     BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_return_output := BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2436_c11_299c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2440_l2433_l2436_DUPLICATE_7f8b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2440_l2433_l2436_DUPLICATE_7f8b_return_output := result.is_stack_write;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2420_c2_fc3f] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2420_c2_fc3f_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2420_c6_fee1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_left;
     BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_return_output := BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2433_l2448_DUPLICATE_4c62 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2433_l2448_DUPLICATE_4c62_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2448_l2436_DUPLICATE_28e9 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2448_l2436_DUPLICATE_28e9_return_output := result.stack_address_sp_offset;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2420_c2_fc3f] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2420_c2_fc3f_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2440_l2433_l2436_DUPLICATE_27db LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2440_l2433_l2436_DUPLICATE_27db_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2440_l2433_l2448_l2436_DUPLICATE_87de LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2440_l2433_l2448_l2436_DUPLICATE_87de_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2420_l2433_l2448_l2436_DUPLICATE_a81a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2420_l2433_l2448_l2436_DUPLICATE_a81a_return_output := result.u8_value;

     -- sp_relative_shift[uxn_opcodes_h_l2438_c30_3f27] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_ins;
     sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_x;
     sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_return_output := sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2433_c11_1b72] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_left;
     BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_return_output := BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2448_c11_184a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2448_c11_184a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c11_184a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2448_c11_184a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c11_184a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c11_184a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2448_c11_184a_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2420_c2_fc3f] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2420_c2_fc3f_return_output := result.is_pc_updated;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c6_fee1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_1b72_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c11_299c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2440_c11_ea1d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c11_184a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c11_184a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c11_184a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2448_c11_184a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2433_l2448_DUPLICATE_4c62_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2433_l2448_DUPLICATE_4c62_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2440_l2433_l2448_l2436_DUPLICATE_87de_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2440_l2433_l2448_l2436_DUPLICATE_87de_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2440_l2433_l2448_l2436_DUPLICATE_87de_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2440_l2433_l2448_l2436_DUPLICATE_87de_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2440_l2433_l2436_DUPLICATE_27db_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2440_l2433_l2436_DUPLICATE_27db_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2440_l2433_l2436_DUPLICATE_27db_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2440_l2433_l2436_DUPLICATE_7f8b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2440_l2433_l2436_DUPLICATE_7f8b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2440_l2433_l2436_DUPLICATE_7f8b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2448_l2436_DUPLICATE_28e9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2448_l2436_DUPLICATE_28e9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2420_l2433_l2448_l2436_DUPLICATE_a81a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2420_l2433_l2448_l2436_DUPLICATE_a81a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2420_l2433_l2448_l2436_DUPLICATE_a81a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2420_l2433_l2448_l2436_DUPLICATE_a81a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2420_c2_fc3f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2420_c2_fc3f_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2420_c2_fc3f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2438_c30_3f27_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2448_c7_decb] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_return_output := result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2448_c7_decb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2440_c7_fedf] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_cond;
     t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output := t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2420_c2_fc3f] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2440_c7_fedf] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2436_c7_07dd] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_cond;
     t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output := t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2440_c7_fedf] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2448_c7_decb] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2448_c7_decb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2420_c2_fc3f] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2420_c2_fc3f] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2448_c7_decb_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2448_c7_decb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2448_c7_decb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2448_c7_decb_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2436_c7_07dd] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2440_c7_fedf] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2440_c7_fedf] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2433_c7_fcec] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_cond;
     t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output := t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2440_c7_fedf] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2440_c7_fedf] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output := result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2436_c7_07dd] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_cond;
     t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output := t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2436_c7_07dd] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2440_c7_fedf_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output;
     -- t16_high_MUX[uxn_opcodes_h_l2420_c2_fc3f] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond;
     t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output := t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2433_c7_fcec] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2433_c7_fcec] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_cond;
     t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output := t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2436_c7_07dd] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output := result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2436_c7_07dd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2433_c7_fcec] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2436_c7_07dd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2436_c7_07dd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2436_c7_07dd_return_output;
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2433_c7_fcec] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2420_c2_fc3f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2433_c7_fcec] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2420_c2_fc3f] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond;
     t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output := t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2433_c7_fcec] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output := result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2433_c7_fcec] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2420_c2_fc3f] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2433_c7_fcec_return_output;
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2420_c2_fc3f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2420_c2_fc3f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2420_c2_fc3f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2420_c2_fc3f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2455_l2416_DUPLICATE_84a1 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2455_l2416_DUPLICATE_84a1_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_04b4(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2420_c2_fc3f_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2455_l2416_DUPLICATE_84a1_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2455_l2416_DUPLICATE_84a1_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
