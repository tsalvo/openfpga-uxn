-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 53
entity ovr_0CLK_6d7675a8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ovr_0CLK_6d7675a8;
architecture arch of ovr_0CLK_6d7675a8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l288_c6_3178]
signal BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l288_c1_11e5]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l288_c2_5632]
signal t8_MUX_uxn_opcodes_h_l288_c2_5632_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l288_c2_5632_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l288_c2_5632_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l288_c2_5632_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l288_c2_5632]
signal result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l288_c2_5632]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l288_c2_5632]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l288_c2_5632]
signal result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l288_c2_5632]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l288_c2_5632]
signal result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l288_c2_5632]
signal n8_MUX_uxn_opcodes_h_l288_c2_5632_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l288_c2_5632_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l288_c2_5632_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l288_c2_5632_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l289_c3_cd8d[uxn_opcodes_h_l289_c3_cd8d]
signal printf_uxn_opcodes_h_l289_c3_cd8d_uxn_opcodes_h_l289_c3_cd8d_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l293_c11_894e]
signal BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l293_c7_664a]
signal t8_MUX_uxn_opcodes_h_l293_c7_664a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l293_c7_664a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l293_c7_664a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l293_c7_664a_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l293_c7_664a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l293_c7_664a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l293_c7_664a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l293_c7_664a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l293_c7_664a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l293_c7_664a]
signal result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l293_c7_664a]
signal n8_MUX_uxn_opcodes_h_l293_c7_664a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l293_c7_664a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l293_c7_664a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l293_c7_664a_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l296_c11_3b45]
signal BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l296_c7_4f37]
signal t8_MUX_uxn_opcodes_h_l296_c7_4f37_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l296_c7_4f37_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l296_c7_4f37]
signal result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l296_c7_4f37]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l296_c7_4f37]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l296_c7_4f37]
signal result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l296_c7_4f37]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l296_c7_4f37]
signal result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l296_c7_4f37]
signal n8_MUX_uxn_opcodes_h_l296_c7_4f37_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l296_c7_4f37_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l299_c11_18e6]
signal BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l299_c7_644d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l299_c7_644d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l299_c7_644d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l299_c7_644d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l299_c7_644d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l299_c7_644d]
signal result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l299_c7_644d]
signal n8_MUX_uxn_opcodes_h_l299_c7_644d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l299_c7_644d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l299_c7_644d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l299_c7_644d_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l302_c30_8963]
signal sp_relative_shift_uxn_opcodes_h_l302_c30_8963_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l302_c30_8963_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l302_c30_8963_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l302_c30_8963_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l307_c11_725b]
signal BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l307_c7_9291]
signal result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l307_c7_9291]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l307_c7_9291]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l307_c7_9291]
signal result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l307_c7_9291]
signal result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l312_c11_c8ee]
signal BIN_OP_EQ_uxn_opcodes_h_l312_c11_c8ee_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l312_c11_c8ee_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l312_c11_c8ee_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l312_c7_ea05]
signal result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l312_c7_ea05]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l312_c7_ea05]
signal result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l312_c7_ea05]
signal result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l316_c11_ab7a]
signal BIN_OP_EQ_uxn_opcodes_h_l316_c11_ab7a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l316_c11_ab7a_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l316_c11_ab7a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l316_c7_2664]
signal result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l316_c7_2664]
signal result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8c29( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178
BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_left,
BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_right,
BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_return_output);

-- t8_MUX_uxn_opcodes_h_l288_c2_5632
t8_MUX_uxn_opcodes_h_l288_c2_5632 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l288_c2_5632_cond,
t8_MUX_uxn_opcodes_h_l288_c2_5632_iftrue,
t8_MUX_uxn_opcodes_h_l288_c2_5632_iffalse,
t8_MUX_uxn_opcodes_h_l288_c2_5632_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632
result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632
result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632
result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632
result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632
result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_cond,
result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_return_output);

-- n8_MUX_uxn_opcodes_h_l288_c2_5632
n8_MUX_uxn_opcodes_h_l288_c2_5632 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l288_c2_5632_cond,
n8_MUX_uxn_opcodes_h_l288_c2_5632_iftrue,
n8_MUX_uxn_opcodes_h_l288_c2_5632_iffalse,
n8_MUX_uxn_opcodes_h_l288_c2_5632_return_output);

-- printf_uxn_opcodes_h_l289_c3_cd8d_uxn_opcodes_h_l289_c3_cd8d
printf_uxn_opcodes_h_l289_c3_cd8d_uxn_opcodes_h_l289_c3_cd8d : entity work.printf_uxn_opcodes_h_l289_c3_cd8d_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l289_c3_cd8d_uxn_opcodes_h_l289_c3_cd8d_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e
BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_left,
BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_right,
BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_return_output);

-- t8_MUX_uxn_opcodes_h_l293_c7_664a
t8_MUX_uxn_opcodes_h_l293_c7_664a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l293_c7_664a_cond,
t8_MUX_uxn_opcodes_h_l293_c7_664a_iftrue,
t8_MUX_uxn_opcodes_h_l293_c7_664a_iffalse,
t8_MUX_uxn_opcodes_h_l293_c7_664a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a
result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a
result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a
result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a
result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a
result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_cond,
result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_return_output);

-- n8_MUX_uxn_opcodes_h_l293_c7_664a
n8_MUX_uxn_opcodes_h_l293_c7_664a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l293_c7_664a_cond,
n8_MUX_uxn_opcodes_h_l293_c7_664a_iftrue,
n8_MUX_uxn_opcodes_h_l293_c7_664a_iffalse,
n8_MUX_uxn_opcodes_h_l293_c7_664a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45
BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_left,
BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_right,
BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_return_output);

-- t8_MUX_uxn_opcodes_h_l296_c7_4f37
t8_MUX_uxn_opcodes_h_l296_c7_4f37 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l296_c7_4f37_cond,
t8_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue,
t8_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse,
t8_MUX_uxn_opcodes_h_l296_c7_4f37_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37
result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37
result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37
result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37
result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37
result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_cond,
result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_return_output);

-- n8_MUX_uxn_opcodes_h_l296_c7_4f37
n8_MUX_uxn_opcodes_h_l296_c7_4f37 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l296_c7_4f37_cond,
n8_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue,
n8_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse,
n8_MUX_uxn_opcodes_h_l296_c7_4f37_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6
BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_left,
BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_right,
BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d
result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d
result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d
result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d
result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d
result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_cond,
result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_return_output);

-- n8_MUX_uxn_opcodes_h_l299_c7_644d
n8_MUX_uxn_opcodes_h_l299_c7_644d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l299_c7_644d_cond,
n8_MUX_uxn_opcodes_h_l299_c7_644d_iftrue,
n8_MUX_uxn_opcodes_h_l299_c7_644d_iffalse,
n8_MUX_uxn_opcodes_h_l299_c7_644d_return_output);

-- sp_relative_shift_uxn_opcodes_h_l302_c30_8963
sp_relative_shift_uxn_opcodes_h_l302_c30_8963 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l302_c30_8963_ins,
sp_relative_shift_uxn_opcodes_h_l302_c30_8963_x,
sp_relative_shift_uxn_opcodes_h_l302_c30_8963_y,
sp_relative_shift_uxn_opcodes_h_l302_c30_8963_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b
BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b_left,
BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b_right,
BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291
result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291
result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_cond,
result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l312_c11_c8ee
BIN_OP_EQ_uxn_opcodes_h_l312_c11_c8ee : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l312_c11_c8ee_left,
BIN_OP_EQ_uxn_opcodes_h_l312_c11_c8ee_right,
BIN_OP_EQ_uxn_opcodes_h_l312_c11_c8ee_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05
result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_cond,
result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l316_c11_ab7a
BIN_OP_EQ_uxn_opcodes_h_l316_c11_ab7a : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l316_c11_ab7a_left,
BIN_OP_EQ_uxn_opcodes_h_l316_c11_ab7a_right,
BIN_OP_EQ_uxn_opcodes_h_l316_c11_ab7a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664
result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664
result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_return_output,
 t8_MUX_uxn_opcodes_h_l288_c2_5632_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_return_output,
 n8_MUX_uxn_opcodes_h_l288_c2_5632_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_return_output,
 t8_MUX_uxn_opcodes_h_l293_c7_664a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_return_output,
 n8_MUX_uxn_opcodes_h_l293_c7_664a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_return_output,
 t8_MUX_uxn_opcodes_h_l296_c7_4f37_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_return_output,
 n8_MUX_uxn_opcodes_h_l296_c7_4f37_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_return_output,
 n8_MUX_uxn_opcodes_h_l299_c7_644d_return_output,
 sp_relative_shift_uxn_opcodes_h_l302_c30_8963_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l312_c11_c8ee_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l316_c11_ab7a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l288_c2_5632_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l288_c2_5632_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l293_c7_664a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l288_c2_5632_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l288_c2_5632_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l290_c3_4a70 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l288_c2_5632_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l288_c2_5632_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l293_c7_664a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l288_c2_5632_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l288_c2_5632_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l289_c3_cd8d_uxn_opcodes_h_l289_c3_cd8d_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l293_c7_664a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l293_c7_664a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l296_c7_4f37_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l293_c7_664a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l294_c3_0b95 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l293_c7_664a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l293_c7_664a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l296_c7_4f37_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l293_c7_664a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l296_c7_4f37_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l299_c7_644d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l296_c7_4f37_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l304_c3_3a7d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l299_c7_644d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l299_c7_644d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l299_c7_644d_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_8963_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_8963_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_8963_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_8963_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l309_c3_ffe8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_c8ee_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_c8ee_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_c8ee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l313_c3_1260 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_ab7a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_ab7a_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_ab7a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l293_l307_l296_l288_DUPLICATE_8bc9_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l316_l312_l307_l296_l293_l288_DUPLICATE_1845_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l293_l296_l288_l299_DUPLICATE_e36d_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l293_l296_l312_l288_DUPLICATE_3cda_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l316_l312_l307_l299_l296_l293_DUPLICATE_9705_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l296_l312_DUPLICATE_8c8e_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l321_l284_DUPLICATE_8b3e_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_c8ee_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_iffalse := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_8963_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l294_c3_0b95 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l294_c3_0b95;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l290_c3_4a70 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l290_c3_4a70;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_ab7a_right := to_unsigned(6, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_8963_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l313_c3_1260 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l313_c3_1260;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l304_c3_3a7d := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l304_c3_3a7d;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l309_c3_ffe8 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l309_c3_ffe8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_8963_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l288_c2_5632_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l293_c7_664a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l299_c7_644d_iffalse := n8;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_iftrue := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_c8ee_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_ab7a_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l299_c7_644d_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l288_c2_5632_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l293_c7_664a_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l299_c11_18e6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_left;
     BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_return_output := BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l296_c11_3b45] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_left;
     BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_return_output := BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l293_l296_l288_l299_DUPLICATE_e36d LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l293_l296_l288_l299_DUPLICATE_e36d_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l307_c11_725b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b_left;
     BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b_return_output := BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l312_c11_c8ee] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l312_c11_c8ee_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_c8ee_left;
     BIN_OP_EQ_uxn_opcodes_h_l312_c11_c8ee_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_c8ee_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_c8ee_return_output := BIN_OP_EQ_uxn_opcodes_h_l312_c11_c8ee_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l293_c11_894e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_left;
     BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_return_output := BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l293_l307_l296_l288_DUPLICATE_8bc9 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l293_l307_l296_l288_DUPLICATE_8bc9_return_output := result.is_sp_shift;

     -- sp_relative_shift[uxn_opcodes_h_l302_c30_8963] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l302_c30_8963_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_8963_ins;
     sp_relative_shift_uxn_opcodes_h_l302_c30_8963_x <= VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_8963_x;
     sp_relative_shift_uxn_opcodes_h_l302_c30_8963_y <= VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_8963_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_8963_return_output := sp_relative_shift_uxn_opcodes_h_l302_c30_8963_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l316_l312_l307_l299_l296_l293_DUPLICATE_9705 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l316_l312_l307_l299_l296_l293_DUPLICATE_9705_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l296_l312_DUPLICATE_8c8e LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l296_l312_DUPLICATE_8c8e_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l316_c11_ab7a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l316_c11_ab7a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_ab7a_left;
     BIN_OP_EQ_uxn_opcodes_h_l316_c11_ab7a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_ab7a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_ab7a_return_output := BIN_OP_EQ_uxn_opcodes_h_l316_c11_ab7a_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l293_l296_l312_l288_DUPLICATE_3cda LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l293_l296_l312_l288_DUPLICATE_3cda_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l316_l312_l307_l296_l293_l288_DUPLICATE_1845 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l316_l312_l307_l296_l293_l288_DUPLICATE_1845_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l288_c6_3178] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_left;
     BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_return_output := BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l288_c2_5632_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l288_c2_5632_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l288_c6_3178_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l293_c7_664a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l293_c7_664a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l293_c11_894e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l296_c7_4f37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l296_c7_4f37_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l296_c11_3b45_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l299_c7_644d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l299_c11_18e6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_725b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_c8ee_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_c8ee_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_c8ee_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l312_c11_c8ee_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_ab7a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l316_c11_ab7a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l293_l296_l288_l299_DUPLICATE_e36d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l293_l296_l288_l299_DUPLICATE_e36d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l293_l296_l288_l299_DUPLICATE_e36d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l293_l296_l288_l299_DUPLICATE_e36d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l316_l312_l307_l299_l296_l293_DUPLICATE_9705_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l316_l312_l307_l299_l296_l293_DUPLICATE_9705_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l316_l312_l307_l299_l296_l293_DUPLICATE_9705_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l316_l312_l307_l299_l296_l293_DUPLICATE_9705_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l316_l312_l307_l299_l296_l293_DUPLICATE_9705_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l316_l312_l307_l299_l296_l293_DUPLICATE_9705_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l293_l307_l296_l288_DUPLICATE_8bc9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l293_l307_l296_l288_DUPLICATE_8bc9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l293_l307_l296_l288_DUPLICATE_8bc9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l293_l307_l296_l288_DUPLICATE_8bc9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l316_l312_l307_l296_l293_l288_DUPLICATE_1845_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l316_l312_l307_l296_l293_l288_DUPLICATE_1845_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l316_l312_l307_l296_l293_l288_DUPLICATE_1845_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l316_l312_l307_l296_l293_l288_DUPLICATE_1845_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l316_l312_l307_l296_l293_l288_DUPLICATE_1845_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l316_l312_l307_l296_l293_l288_DUPLICATE_1845_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l296_l312_DUPLICATE_8c8e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l296_l312_DUPLICATE_8c8e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l293_l296_l312_l288_DUPLICATE_3cda_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l293_l296_l312_l288_DUPLICATE_3cda_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l293_l296_l312_l288_DUPLICATE_3cda_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l293_l296_l312_l288_DUPLICATE_3cda_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l302_c30_8963_return_output;
     -- t8_MUX[uxn_opcodes_h_l296_c7_4f37] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l296_c7_4f37_cond <= VAR_t8_MUX_uxn_opcodes_h_l296_c7_4f37_cond;
     t8_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue;
     t8_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l296_c7_4f37_return_output := t8_MUX_uxn_opcodes_h_l296_c7_4f37_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l316_c7_2664] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l307_c7_9291] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l312_c7_ea05] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l288_c1_11e5] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l316_c7_2664] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_return_output;

     -- n8_MUX[uxn_opcodes_h_l299_c7_644d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l299_c7_644d_cond <= VAR_n8_MUX_uxn_opcodes_h_l299_c7_644d_cond;
     n8_MUX_uxn_opcodes_h_l299_c7_644d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l299_c7_644d_iftrue;
     n8_MUX_uxn_opcodes_h_l299_c7_644d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l299_c7_644d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l299_c7_644d_return_output := n8_MUX_uxn_opcodes_h_l299_c7_644d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l299_c7_644d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l312_c7_ea05] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_cond;
     result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_return_output := result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l289_c3_cd8d_uxn_opcodes_h_l289_c3_cd8d_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l288_c1_11e5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse := VAR_n8_MUX_uxn_opcodes_h_l299_c7_644d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l316_c7_2664_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l307_c7_9291_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l316_c7_2664_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l299_c7_644d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l312_c7_ea05_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l312_c7_ea05_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l293_c7_664a_iffalse := VAR_t8_MUX_uxn_opcodes_h_l296_c7_4f37_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l307_c7_9291] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l307_c7_9291] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_cond;
     result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_return_output := result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l299_c7_644d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l312_c7_ea05] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_return_output;

     -- t8_MUX[uxn_opcodes_h_l293_c7_664a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l293_c7_664a_cond <= VAR_t8_MUX_uxn_opcodes_h_l293_c7_664a_cond;
     t8_MUX_uxn_opcodes_h_l293_c7_664a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l293_c7_664a_iftrue;
     t8_MUX_uxn_opcodes_h_l293_c7_664a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l293_c7_664a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l293_c7_664a_return_output := t8_MUX_uxn_opcodes_h_l293_c7_664a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l312_c7_ea05] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_return_output;

     -- n8_MUX[uxn_opcodes_h_l296_c7_4f37] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l296_c7_4f37_cond <= VAR_n8_MUX_uxn_opcodes_h_l296_c7_4f37_cond;
     n8_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue;
     n8_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l296_c7_4f37_return_output := n8_MUX_uxn_opcodes_h_l296_c7_4f37_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l296_c7_4f37] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_return_output;

     -- printf_uxn_opcodes_h_l289_c3_cd8d[uxn_opcodes_h_l289_c3_cd8d] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l289_c3_cd8d_uxn_opcodes_h_l289_c3_cd8d_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l289_c3_cd8d_uxn_opcodes_h_l289_c3_cd8d_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l293_c7_664a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l296_c7_4f37_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l312_c7_ea05_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l299_c7_644d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l312_c7_ea05_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l296_c7_4f37_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_9291_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_9291_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l288_c2_5632_iffalse := VAR_t8_MUX_uxn_opcodes_h_l293_c7_664a_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l307_c7_9291] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l307_c7_9291] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_return_output;

     -- n8_MUX[uxn_opcodes_h_l293_c7_664a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l293_c7_664a_cond <= VAR_n8_MUX_uxn_opcodes_h_l293_c7_664a_cond;
     n8_MUX_uxn_opcodes_h_l293_c7_664a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l293_c7_664a_iftrue;
     n8_MUX_uxn_opcodes_h_l293_c7_664a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l293_c7_664a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l293_c7_664a_return_output := n8_MUX_uxn_opcodes_h_l293_c7_664a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l293_c7_664a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l299_c7_644d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_return_output;

     -- t8_MUX[uxn_opcodes_h_l288_c2_5632] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l288_c2_5632_cond <= VAR_t8_MUX_uxn_opcodes_h_l288_c2_5632_cond;
     t8_MUX_uxn_opcodes_h_l288_c2_5632_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l288_c2_5632_iftrue;
     t8_MUX_uxn_opcodes_h_l288_c2_5632_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l288_c2_5632_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l288_c2_5632_return_output := t8_MUX_uxn_opcodes_h_l288_c2_5632_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l299_c7_644d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_return_output := result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l296_c7_4f37] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l288_c2_5632_iffalse := VAR_n8_MUX_uxn_opcodes_h_l293_c7_664a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_9291_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l296_c7_4f37_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_9291_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l293_c7_664a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l299_c7_644d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l299_c7_644d_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l288_c2_5632_return_output;
     -- n8_MUX[uxn_opcodes_h_l288_c2_5632] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l288_c2_5632_cond <= VAR_n8_MUX_uxn_opcodes_h_l288_c2_5632_cond;
     n8_MUX_uxn_opcodes_h_l288_c2_5632_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l288_c2_5632_iftrue;
     n8_MUX_uxn_opcodes_h_l288_c2_5632_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l288_c2_5632_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l288_c2_5632_return_output := n8_MUX_uxn_opcodes_h_l288_c2_5632_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l299_c7_644d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l293_c7_664a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l296_c7_4f37] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_cond;
     result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_return_output := result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l299_c7_644d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l288_c2_5632] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l296_c7_4f37] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l288_c2_5632_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l299_c7_644d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l293_c7_664a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l299_c7_644d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l296_c7_4f37_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l296_c7_4f37_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l288_c2_5632] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l293_c7_664a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l293_c7_664a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_return_output := result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l296_c7_4f37] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l296_c7_4f37] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l296_c7_4f37_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l296_c7_4f37_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l293_c7_664a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l293_c7_664a_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l288_c2_5632] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l293_c7_664a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l293_c7_664a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l288_c2_5632] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_cond;
     result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_return_output := result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_return_output;

     -- Submodule level 7
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l293_c7_664a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l293_c7_664a_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l288_c2_5632] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l288_c2_5632] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_return_output;

     -- Submodule level 8
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l321_l284_DUPLICATE_8b3e LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l321_l284_DUPLICATE_8b3e_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8c29(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l288_c2_5632_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l288_c2_5632_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l288_c2_5632_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l288_c2_5632_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l288_c2_5632_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l288_c2_5632_return_output);

     -- Submodule level 9
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l321_l284_DUPLICATE_8b3e_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l321_l284_DUPLICATE_8b3e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
