-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 80
entity deo2_0CLK_41131849 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_device_ram_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end deo2_0CLK_41131849;
architecture arch of deo2_0CLK_41131849 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal l8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal current_deo_phase : unsigned(7 downto 0) := to_unsigned(0, 8);
signal deo_param0 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal deo_param1 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal is_second_deo : unsigned(0 downto 0) := to_unsigned(0, 1);
signal is_phase_3 : unsigned(0 downto 0) := to_unsigned(0, 1);
signal is_phase_4 : unsigned(0 downto 0) := to_unsigned(0, 1);
signal result : opcode_result_t := opcode_result_t_NULL;
signal device_out_result : device_out_result_t := device_out_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_l8 : unsigned(7 downto 0);
signal REG_COMB_current_deo_phase : unsigned(7 downto 0);
signal REG_COMB_deo_param0 : unsigned(7 downto 0);
signal REG_COMB_deo_param1 : unsigned(7 downto 0);
signal REG_COMB_is_second_deo : unsigned(0 downto 0);
signal REG_COMB_is_phase_3 : unsigned(0 downto 0);
signal REG_COMB_is_phase_4 : unsigned(0 downto 0);
signal REG_COMB_result : opcode_result_t;
signal REG_COMB_device_out_result : device_out_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l539_c6_9f48]
signal BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l548_c7_ce40]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(0 downto 0);

-- is_phase_4_MUX[uxn_opcodes_h_l539_c2_8124]
signal is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
signal is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(0 downto 0);
signal is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(0 downto 0);
signal is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l539_c2_8124]
signal l8_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l539_c2_8124]
signal result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(7 downto 0);

-- result_vram_write_layer_MUX[uxn_opcodes_h_l539_c2_8124]
signal result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l539_c2_8124]
signal result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l539_c2_8124]
signal result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(15 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l539_c2_8124]
signal result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l539_c2_8124]
signal result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(0 downto 0);

-- result_is_device_ram_write_MUX[uxn_opcodes_h_l539_c2_8124]
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l539_c2_8124]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l539_c2_8124]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(3 downto 0);

-- is_second_deo_MUX[uxn_opcodes_h_l539_c2_8124]
signal is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(0 downto 0);

-- current_deo_phase_MUX[uxn_opcodes_h_l539_c2_8124]
signal current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(7 downto 0);

-- deo_param1_MUX[uxn_opcodes_h_l539_c2_8124]
signal deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(7 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(7 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(7 downto 0);

-- device_out_result_MUX[uxn_opcodes_h_l539_c2_8124]
signal device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
signal device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_return_output : device_out_result_t;

-- deo_param0_MUX[uxn_opcodes_h_l539_c2_8124]
signal deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(7 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(7 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l539_c2_8124]
signal n8_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(7 downto 0);

-- is_phase_3_MUX[uxn_opcodes_h_l539_c2_8124]
signal is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
signal is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(0 downto 0);
signal is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(0 downto 0);
signal is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l539_c2_8124]
signal t8_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l548_c11_6174]
signal BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l551_c7_205d]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(0 downto 0);

-- is_phase_4_MUX[uxn_opcodes_h_l548_c7_ce40]
signal is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
signal is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(0 downto 0);
signal is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(0 downto 0);
signal is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l548_c7_ce40]
signal l8_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l548_c7_ce40]
signal result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(7 downto 0);

-- result_vram_write_layer_MUX[uxn_opcodes_h_l548_c7_ce40]
signal result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l548_c7_ce40]
signal result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l548_c7_ce40]
signal result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(15 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l548_c7_ce40]
signal result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l548_c7_ce40]
signal result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(0 downto 0);

-- result_is_device_ram_write_MUX[uxn_opcodes_h_l548_c7_ce40]
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l548_c7_ce40]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l548_c7_ce40]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(3 downto 0);

-- is_second_deo_MUX[uxn_opcodes_h_l548_c7_ce40]
signal is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(0 downto 0);

-- current_deo_phase_MUX[uxn_opcodes_h_l548_c7_ce40]
signal current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(7 downto 0);

-- deo_param1_MUX[uxn_opcodes_h_l548_c7_ce40]
signal deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(7 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(7 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(7 downto 0);

-- device_out_result_MUX[uxn_opcodes_h_l548_c7_ce40]
signal device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
signal device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : device_out_result_t;

-- deo_param0_MUX[uxn_opcodes_h_l548_c7_ce40]
signal deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(7 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(7 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l548_c7_ce40]
signal n8_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(7 downto 0);

-- is_phase_3_MUX[uxn_opcodes_h_l548_c7_ce40]
signal is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
signal is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(0 downto 0);
signal is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(0 downto 0);
signal is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l548_c7_ce40]
signal t8_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l551_c11_ffc2]
signal BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l555_c1_b0c5]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_return_output : unsigned(0 downto 0);

-- is_phase_4_MUX[uxn_opcodes_h_l551_c7_205d]
signal is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
signal is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(0 downto 0);
signal is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(0 downto 0);
signal is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l551_c7_205d]
signal l8_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l551_c7_205d]
signal result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(7 downto 0);

-- result_vram_write_layer_MUX[uxn_opcodes_h_l551_c7_205d]
signal result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l551_c7_205d]
signal result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l551_c7_205d]
signal result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(15 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l551_c7_205d]
signal result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l551_c7_205d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(0 downto 0);

-- result_is_device_ram_write_MUX[uxn_opcodes_h_l551_c7_205d]
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l551_c7_205d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l551_c7_205d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(3 downto 0);

-- is_second_deo_MUX[uxn_opcodes_h_l551_c7_205d]
signal is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(0 downto 0);

-- current_deo_phase_MUX[uxn_opcodes_h_l551_c7_205d]
signal current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(7 downto 0);

-- deo_param1_MUX[uxn_opcodes_h_l551_c7_205d]
signal deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(7 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(7 downto 0);
signal deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(7 downto 0);

-- device_out_result_MUX[uxn_opcodes_h_l551_c7_205d]
signal device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
signal device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_return_output : device_out_result_t;

-- deo_param0_MUX[uxn_opcodes_h_l551_c7_205d]
signal deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(7 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(7 downto 0);
signal deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l551_c7_205d]
signal n8_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(7 downto 0);

-- is_phase_3_MUX[uxn_opcodes_h_l551_c7_205d]
signal is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
signal is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(0 downto 0);
signal is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(0 downto 0);
signal is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l551_c7_205d]
signal t8_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l556_c17_5fcc]
signal BIN_OP_EQ_uxn_opcodes_h_l556_c17_5fcc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l556_c17_5fcc_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l556_c17_5fcc_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l556_c17_aaf6]
signal MUX_uxn_opcodes_h_l556_c17_aaf6_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l556_c17_aaf6_iftrue : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l556_c17_aaf6_iffalse : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l556_c17_aaf6_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l557_c17_c8c7]
signal BIN_OP_EQ_uxn_opcodes_h_l557_c17_c8c7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l557_c17_c8c7_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l557_c17_c8c7_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l557_c17_bfc8]
signal MUX_uxn_opcodes_h_l557_c17_bfc8_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l557_c17_bfc8_iftrue : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l557_c17_bfc8_iffalse : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l557_c17_bfc8_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l558_c8_9c1c]
signal MUX_uxn_opcodes_h_l558_c8_9c1c_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l558_c8_9c1c_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l558_c8_9c1c_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l558_c8_9c1c_return_output : unsigned(7 downto 0);

-- MUX[uxn_opcodes_h_l559_c8_9d6a]
signal MUX_uxn_opcodes_h_l559_c8_9d6a_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l559_c8_9d6a_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l559_c8_9d6a_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l559_c8_9d6a_return_output : unsigned(7 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l560_c32_60a0]
signal BIN_OP_PLUS_uxn_opcodes_h_l560_c32_60a0_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l560_c32_60a0_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l560_c32_60a0_return_output : unsigned(8 downto 0);

-- MUX[uxn_opcodes_h_l560_c16_ee8b]
signal MUX_uxn_opcodes_h_l560_c16_ee8b_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l560_c16_ee8b_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l560_c16_ee8b_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l560_c16_ee8b_return_output : unsigned(7 downto 0);

-- MUX[uxn_opcodes_h_l561_c16_e93e]
signal MUX_uxn_opcodes_h_l561_c16_e93e_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l561_c16_e93e_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l561_c16_e93e_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l561_c16_e93e_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l562_c43_1dbf]
signal sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_return_output : signed(3 downto 0);

-- MUX[uxn_opcodes_h_l562_c30_d095]
signal MUX_uxn_opcodes_h_l562_c30_d095_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l562_c30_d095_iftrue : signed(3 downto 0);
signal MUX_uxn_opcodes_h_l562_c30_d095_iffalse : signed(3 downto 0);
signal MUX_uxn_opcodes_h_l562_c30_d095_return_output : signed(3 downto 0);

-- device_out[uxn_opcodes_h_l563_c23_d468]
signal device_out_uxn_opcodes_h_l563_c23_d468_CLOCK_ENABLE : unsigned(0 downto 0);
signal device_out_uxn_opcodes_h_l563_c23_d468_device_address : unsigned(7 downto 0);
signal device_out_uxn_opcodes_h_l563_c23_d468_value : unsigned(7 downto 0);
signal device_out_uxn_opcodes_h_l563_c23_d468_phase : unsigned(7 downto 0);
signal device_out_uxn_opcodes_h_l563_c23_d468_previous_device_ram_read : unsigned(7 downto 0);
signal device_out_uxn_opcodes_h_l563_c23_d468_previous_ram_read : unsigned(7 downto 0);
signal device_out_uxn_opcodes_h_l563_c23_d468_return_output : device_out_result_t;

-- BIN_OP_AND[uxn_opcodes_h_l570_c24_c405]
signal BIN_OP_AND_uxn_opcodes_h_l570_c24_c405_left : unsigned(0 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l570_c24_c405_right : unsigned(0 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l570_c24_c405_return_output : unsigned(0 downto 0);

-- is_second_deo_MUX[uxn_opcodes_h_l571_c3_6837]
signal is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_cond : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_iftrue : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_iffalse : unsigned(0 downto 0);
signal is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_return_output : unsigned(0 downto 0);

-- current_deo_phase_MUX[uxn_opcodes_h_l571_c3_6837]
signal current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_cond : unsigned(0 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_iftrue : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_iffalse : unsigned(7 downto 0);
signal current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_return_output : unsigned(7 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l575_c4_0ea3]
signal BIN_OP_PLUS_uxn_opcodes_h_l575_c4_0ea3_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l575_c4_0ea3_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l575_c4_0ea3_return_output : unsigned(8 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_f18e( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : signed;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.vram_write_layer := ref_toks_2;
      base.is_vram_write := ref_toks_3;
      base.u16_value := ref_toks_4;
      base.device_ram_address := ref_toks_5;
      base.is_opc_done := ref_toks_6;
      base.is_device_ram_write := ref_toks_7;
      base.sp_relative_shift := ref_toks_8;
      base.stack_address_sp_offset := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48
BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_left,
BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_right,
BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_return_output);

-- is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124
is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_cond,
is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_iftrue,
is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_iffalse,
is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_return_output);

-- l8_MUX_uxn_opcodes_h_l539_c2_8124
l8_MUX_uxn_opcodes_h_l539_c2_8124 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l539_c2_8124_cond,
l8_MUX_uxn_opcodes_h_l539_c2_8124_iftrue,
l8_MUX_uxn_opcodes_h_l539_c2_8124_iffalse,
l8_MUX_uxn_opcodes_h_l539_c2_8124_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124
result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_cond,
result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_return_output);

-- result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124
result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_cond,
result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_iftrue,
result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_iffalse,
result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124
result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124
result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_cond,
result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124
result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124
result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_return_output);

-- result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124
result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_cond,
result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_iftrue,
result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_iffalse,
result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124
result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_return_output);

-- is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124
is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_cond,
is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_iftrue,
is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_iffalse,
is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_return_output);

-- current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124
current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_cond,
current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_iftrue,
current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_iffalse,
current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_return_output);

-- deo_param1_MUX_uxn_opcodes_h_l539_c2_8124
deo_param1_MUX_uxn_opcodes_h_l539_c2_8124 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_cond,
deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_iftrue,
deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_iffalse,
deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_return_output);

-- device_out_result_MUX_uxn_opcodes_h_l539_c2_8124
device_out_result_MUX_uxn_opcodes_h_l539_c2_8124 : entity work.MUX_uint1_t_device_out_result_t_device_out_result_t_0CLK_de264c78 port map (
device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_cond,
device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_iftrue,
device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_iffalse,
device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_return_output);

-- deo_param0_MUX_uxn_opcodes_h_l539_c2_8124
deo_param0_MUX_uxn_opcodes_h_l539_c2_8124 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_cond,
deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_iftrue,
deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_iffalse,
deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_return_output);

-- n8_MUX_uxn_opcodes_h_l539_c2_8124
n8_MUX_uxn_opcodes_h_l539_c2_8124 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l539_c2_8124_cond,
n8_MUX_uxn_opcodes_h_l539_c2_8124_iftrue,
n8_MUX_uxn_opcodes_h_l539_c2_8124_iffalse,
n8_MUX_uxn_opcodes_h_l539_c2_8124_return_output);

-- is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124
is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_cond,
is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_iftrue,
is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_iffalse,
is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_return_output);

-- t8_MUX_uxn_opcodes_h_l539_c2_8124
t8_MUX_uxn_opcodes_h_l539_c2_8124 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l539_c2_8124_cond,
t8_MUX_uxn_opcodes_h_l539_c2_8124_iftrue,
t8_MUX_uxn_opcodes_h_l539_c2_8124_iffalse,
t8_MUX_uxn_opcodes_h_l539_c2_8124_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174
BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_left,
BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_right,
BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_return_output);

-- is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40
is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_cond,
is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue,
is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse,
is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_return_output);

-- l8_MUX_uxn_opcodes_h_l548_c7_ce40
l8_MUX_uxn_opcodes_h_l548_c7_ce40 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l548_c7_ce40_cond,
l8_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue,
l8_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse,
l8_MUX_uxn_opcodes_h_l548_c7_ce40_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40
result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_cond,
result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_return_output);

-- result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40
result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_cond,
result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue,
result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse,
result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40
result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40
result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_cond,
result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40
result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40
result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_return_output);

-- result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40
result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_cond,
result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue,
result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse,
result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40
result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_return_output);

-- is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40
is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_cond,
is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue,
is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse,
is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_return_output);

-- current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40
current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_cond,
current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue,
current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse,
current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_return_output);

-- deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40
deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_cond,
deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue,
deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse,
deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_return_output);

-- device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40
device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40 : entity work.MUX_uint1_t_device_out_result_t_device_out_result_t_0CLK_de264c78 port map (
device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_cond,
device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue,
device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse,
device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_return_output);

-- deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40
deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_cond,
deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue,
deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse,
deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_return_output);

-- n8_MUX_uxn_opcodes_h_l548_c7_ce40
n8_MUX_uxn_opcodes_h_l548_c7_ce40 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l548_c7_ce40_cond,
n8_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue,
n8_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse,
n8_MUX_uxn_opcodes_h_l548_c7_ce40_return_output);

-- is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40
is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_cond,
is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue,
is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse,
is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_return_output);

-- t8_MUX_uxn_opcodes_h_l548_c7_ce40
t8_MUX_uxn_opcodes_h_l548_c7_ce40 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l548_c7_ce40_cond,
t8_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue,
t8_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse,
t8_MUX_uxn_opcodes_h_l548_c7_ce40_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2
BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_left,
BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_right,
BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_return_output);

-- is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d
is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_cond,
is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_iftrue,
is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_iffalse,
is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_return_output);

-- l8_MUX_uxn_opcodes_h_l551_c7_205d
l8_MUX_uxn_opcodes_h_l551_c7_205d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l551_c7_205d_cond,
l8_MUX_uxn_opcodes_h_l551_c7_205d_iftrue,
l8_MUX_uxn_opcodes_h_l551_c7_205d_iffalse,
l8_MUX_uxn_opcodes_h_l551_c7_205d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d
result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_cond,
result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_return_output);

-- result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d
result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_cond,
result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_iftrue,
result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_iffalse,
result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d
result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d
result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_cond,
result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d
result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d
result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_return_output);

-- result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d
result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_cond,
result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_iftrue,
result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_iffalse,
result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d
result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_return_output);

-- is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d
is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_cond,
is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_iftrue,
is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_iffalse,
is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_return_output);

-- current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d
current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_cond,
current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_iftrue,
current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_iffalse,
current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_return_output);

-- deo_param1_MUX_uxn_opcodes_h_l551_c7_205d
deo_param1_MUX_uxn_opcodes_h_l551_c7_205d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_cond,
deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_iftrue,
deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_iffalse,
deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_return_output);

-- device_out_result_MUX_uxn_opcodes_h_l551_c7_205d
device_out_result_MUX_uxn_opcodes_h_l551_c7_205d : entity work.MUX_uint1_t_device_out_result_t_device_out_result_t_0CLK_de264c78 port map (
device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_cond,
device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_iftrue,
device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_iffalse,
device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_return_output);

-- deo_param0_MUX_uxn_opcodes_h_l551_c7_205d
deo_param0_MUX_uxn_opcodes_h_l551_c7_205d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_cond,
deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_iftrue,
deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_iffalse,
deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_return_output);

-- n8_MUX_uxn_opcodes_h_l551_c7_205d
n8_MUX_uxn_opcodes_h_l551_c7_205d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l551_c7_205d_cond,
n8_MUX_uxn_opcodes_h_l551_c7_205d_iftrue,
n8_MUX_uxn_opcodes_h_l551_c7_205d_iffalse,
n8_MUX_uxn_opcodes_h_l551_c7_205d_return_output);

-- is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d
is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_cond,
is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_iftrue,
is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_iffalse,
is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_return_output);

-- t8_MUX_uxn_opcodes_h_l551_c7_205d
t8_MUX_uxn_opcodes_h_l551_c7_205d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l551_c7_205d_cond,
t8_MUX_uxn_opcodes_h_l551_c7_205d_iftrue,
t8_MUX_uxn_opcodes_h_l551_c7_205d_iffalse,
t8_MUX_uxn_opcodes_h_l551_c7_205d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l556_c17_5fcc
BIN_OP_EQ_uxn_opcodes_h_l556_c17_5fcc : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l556_c17_5fcc_left,
BIN_OP_EQ_uxn_opcodes_h_l556_c17_5fcc_right,
BIN_OP_EQ_uxn_opcodes_h_l556_c17_5fcc_return_output);

-- MUX_uxn_opcodes_h_l556_c17_aaf6
MUX_uxn_opcodes_h_l556_c17_aaf6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l556_c17_aaf6_cond,
MUX_uxn_opcodes_h_l556_c17_aaf6_iftrue,
MUX_uxn_opcodes_h_l556_c17_aaf6_iffalse,
MUX_uxn_opcodes_h_l556_c17_aaf6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l557_c17_c8c7
BIN_OP_EQ_uxn_opcodes_h_l557_c17_c8c7 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l557_c17_c8c7_left,
BIN_OP_EQ_uxn_opcodes_h_l557_c17_c8c7_right,
BIN_OP_EQ_uxn_opcodes_h_l557_c17_c8c7_return_output);

-- MUX_uxn_opcodes_h_l557_c17_bfc8
MUX_uxn_opcodes_h_l557_c17_bfc8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l557_c17_bfc8_cond,
MUX_uxn_opcodes_h_l557_c17_bfc8_iftrue,
MUX_uxn_opcodes_h_l557_c17_bfc8_iffalse,
MUX_uxn_opcodes_h_l557_c17_bfc8_return_output);

-- MUX_uxn_opcodes_h_l558_c8_9c1c
MUX_uxn_opcodes_h_l558_c8_9c1c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l558_c8_9c1c_cond,
MUX_uxn_opcodes_h_l558_c8_9c1c_iftrue,
MUX_uxn_opcodes_h_l558_c8_9c1c_iffalse,
MUX_uxn_opcodes_h_l558_c8_9c1c_return_output);

-- MUX_uxn_opcodes_h_l559_c8_9d6a
MUX_uxn_opcodes_h_l559_c8_9d6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l559_c8_9d6a_cond,
MUX_uxn_opcodes_h_l559_c8_9d6a_iftrue,
MUX_uxn_opcodes_h_l559_c8_9d6a_iffalse,
MUX_uxn_opcodes_h_l559_c8_9d6a_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l560_c32_60a0
BIN_OP_PLUS_uxn_opcodes_h_l560_c32_60a0 : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l560_c32_60a0_left,
BIN_OP_PLUS_uxn_opcodes_h_l560_c32_60a0_right,
BIN_OP_PLUS_uxn_opcodes_h_l560_c32_60a0_return_output);

-- MUX_uxn_opcodes_h_l560_c16_ee8b
MUX_uxn_opcodes_h_l560_c16_ee8b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l560_c16_ee8b_cond,
MUX_uxn_opcodes_h_l560_c16_ee8b_iftrue,
MUX_uxn_opcodes_h_l560_c16_ee8b_iffalse,
MUX_uxn_opcodes_h_l560_c16_ee8b_return_output);

-- MUX_uxn_opcodes_h_l561_c16_e93e
MUX_uxn_opcodes_h_l561_c16_e93e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l561_c16_e93e_cond,
MUX_uxn_opcodes_h_l561_c16_e93e_iftrue,
MUX_uxn_opcodes_h_l561_c16_e93e_iffalse,
MUX_uxn_opcodes_h_l561_c16_e93e_return_output);

-- sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf
sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_ins,
sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_x,
sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_y,
sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_return_output);

-- MUX_uxn_opcodes_h_l562_c30_d095
MUX_uxn_opcodes_h_l562_c30_d095 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l562_c30_d095_cond,
MUX_uxn_opcodes_h_l562_c30_d095_iftrue,
MUX_uxn_opcodes_h_l562_c30_d095_iffalse,
MUX_uxn_opcodes_h_l562_c30_d095_return_output);

-- device_out_uxn_opcodes_h_l563_c23_d468
device_out_uxn_opcodes_h_l563_c23_d468 : entity work.device_out_0CLK_95124a2a port map (
clk,
device_out_uxn_opcodes_h_l563_c23_d468_CLOCK_ENABLE,
device_out_uxn_opcodes_h_l563_c23_d468_device_address,
device_out_uxn_opcodes_h_l563_c23_d468_value,
device_out_uxn_opcodes_h_l563_c23_d468_phase,
device_out_uxn_opcodes_h_l563_c23_d468_previous_device_ram_read,
device_out_uxn_opcodes_h_l563_c23_d468_previous_ram_read,
device_out_uxn_opcodes_h_l563_c23_d468_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l570_c24_c405
BIN_OP_AND_uxn_opcodes_h_l570_c24_c405 : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l570_c24_c405_left,
BIN_OP_AND_uxn_opcodes_h_l570_c24_c405_right,
BIN_OP_AND_uxn_opcodes_h_l570_c24_c405_return_output);

-- is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837
is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_cond,
is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_iftrue,
is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_iffalse,
is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_return_output);

-- current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837
current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_cond,
current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_iftrue,
current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_iffalse,
current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l575_c4_0ea3
BIN_OP_PLUS_uxn_opcodes_h_l575_c4_0ea3 : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l575_c4_0ea3_left,
BIN_OP_PLUS_uxn_opcodes_h_l575_c4_0ea3_right,
BIN_OP_PLUS_uxn_opcodes_h_l575_c4_0ea3_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_device_ram_read,
 previous_ram_read,
 -- Registers
 t8,
 n8,
 l8,
 current_deo_phase,
 deo_param0,
 deo_param1,
 is_second_deo,
 is_phase_3,
 is_phase_4,
 result,
 device_out_result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_return_output,
 is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
 l8_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
 result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
 result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
 is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
 current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
 deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
 device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
 deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
 n8_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
 is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
 t8_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_return_output,
 is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_return_output,
 l8_MUX_uxn_opcodes_h_l548_c7_ce40_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_return_output,
 result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_return_output,
 result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_return_output,
 is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_return_output,
 current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_return_output,
 deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_return_output,
 device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_return_output,
 deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_return_output,
 n8_MUX_uxn_opcodes_h_l548_c7_ce40_return_output,
 is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_return_output,
 t8_MUX_uxn_opcodes_h_l548_c7_ce40_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_return_output,
 is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_return_output,
 l8_MUX_uxn_opcodes_h_l551_c7_205d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_return_output,
 result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_return_output,
 result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_return_output,
 is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_return_output,
 current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_return_output,
 deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_return_output,
 device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_return_output,
 deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_return_output,
 n8_MUX_uxn_opcodes_h_l551_c7_205d_return_output,
 is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_return_output,
 t8_MUX_uxn_opcodes_h_l551_c7_205d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l556_c17_5fcc_return_output,
 MUX_uxn_opcodes_h_l556_c17_aaf6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l557_c17_c8c7_return_output,
 MUX_uxn_opcodes_h_l557_c17_bfc8_return_output,
 MUX_uxn_opcodes_h_l558_c8_9c1c_return_output,
 MUX_uxn_opcodes_h_l559_c8_9d6a_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l560_c32_60a0_return_output,
 MUX_uxn_opcodes_h_l560_c16_ee8b_return_output,
 MUX_uxn_opcodes_h_l561_c16_e93e_return_output,
 sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_return_output,
 MUX_uxn_opcodes_h_l562_c30_d095_return_output,
 device_out_uxn_opcodes_h_l563_c23_d468_return_output,
 BIN_OP_AND_uxn_opcodes_h_l570_c24_c405_return_output,
 is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_return_output,
 current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l575_c4_0ea3_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(0 downto 0);
 variable VAR_is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(0 downto 0);
 variable VAR_is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(0 downto 0);
 variable VAR_is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(0 downto 0);
 variable VAR_is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(0 downto 0);
 variable VAR_is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l543_c3_51f3 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(7 downto 0);
 variable VAR_current_deo_phase_uxn_opcodes_h_l546_c3_3298 : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_return_output : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
 variable VAR_is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(0 downto 0);
 variable VAR_is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(0 downto 0);
 variable VAR_is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(0 downto 0);
 variable VAR_is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(0 downto 0);
 variable VAR_is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l539_c2_8124_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l539_c2_8124_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l548_c7_ce40_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l539_c2_8124_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l539_c2_8124_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(0 downto 0);
 variable VAR_is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(0 downto 0);
 variable VAR_is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(0 downto 0);
 variable VAR_is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(0 downto 0);
 variable VAR_is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l549_c3_9a1e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_return_output : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
 variable VAR_is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(0 downto 0);
 variable VAR_is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(0 downto 0);
 variable VAR_is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(0 downto 0);
 variable VAR_is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l548_c7_ce40_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_iffalse : unsigned(0 downto 0);
 variable VAR_is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(0 downto 0);
 variable VAR_is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(0 downto 0);
 variable VAR_is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l552_c3_f51c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l551_c7_205d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_return_output : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_return_output : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(7 downto 0);
 variable VAR_deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(7 downto 0);
 variable VAR_deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
 variable VAR_is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(0 downto 0);
 variable VAR_is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(0 downto 0);
 variable VAR_is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l551_c7_205d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l551_c7_205d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l551_c7_205d_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l556_c17_aaf6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c17_5fcc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c17_5fcc_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c17_5fcc_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l556_c17_aaf6_iftrue : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l556_c17_aaf6_iffalse : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l556_c17_aaf6_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l557_c17_bfc8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l557_c17_c8c7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l557_c17_c8c7_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l557_c17_c8c7_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l557_c17_bfc8_iftrue : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l557_c17_bfc8_iffalse : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l557_c17_bfc8_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l558_c8_9c1c_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l558_c8_9c1c_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l558_c8_9c1c_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l558_c8_9c1c_return_output : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l559_c8_9d6a_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l559_c8_9d6a_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l559_c8_9d6a_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l559_c8_9d6a_return_output : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l560_c16_ee8b_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l560_c16_ee8b_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l560_c16_ee8b_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l560_c32_60a0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l560_c32_60a0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l560_c32_60a0_return_output : unsigned(8 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l560_c16_ee8b_return_output : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l561_c16_e93e_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l561_c16_e93e_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l561_c16_e93e_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l561_c16_e93e_return_output : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l562_c30_d095_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l562_c30_d095_iftrue : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l562_c30_d095_iffalse : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l562_c30_d095_return_output : signed(3 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l563_c23_d468_device_address : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l563_c23_d468_value : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l563_c23_d468_phase : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l563_c23_d468_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l563_c23_d468_previous_ram_read : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l563_c23_d468_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l563_c23_d468_return_output : device_out_result_t;
 variable VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l564_c32_f2a0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_device_out_result_t_device_ram_address_d41d_uxn_opcodes_h_l565_c31_6b03_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_vram_write_d41d_uxn_opcodes_h_l566_c26_75a1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_device_out_result_t_vram_write_layer_d41d_uxn_opcodes_h_l567_c29_f9a5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_device_out_result_t_u16_addr_d41d_uxn_opcodes_h_l568_c22_b6cb_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_device_out_result_t_u8_value_d41d_uxn_opcodes_h_l569_c21_f77c_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l570_c24_c405_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l570_c24_c405_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l570_c24_c405_return_output : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_iftrue : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_iffalse : unsigned(0 downto 0);
 variable VAR_is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_cond : unsigned(0 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_iftrue : unsigned(7 downto 0);
 variable VAR_current_deo_phase_uxn_opcodes_h_l572_c4_b061 : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_iffalse : unsigned(7 downto 0);
 variable VAR_current_deo_phase_uxn_opcodes_h_l575_c4_f6a7 : unsigned(7 downto 0);
 variable VAR_current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l575_c4_0ea3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l575_c4_0ea3_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l575_c4_0ea3_return_output : unsigned(8 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_4e2e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_176c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_c949_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_127b_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_8fa6_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_271a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_85a2_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l548_l551_DUPLICATE_336e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d_uxn_opcodes_h_l570_l571_DUPLICATE_f81b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_f18e_uxn_opcodes_h_l579_l533_DUPLICATE_d422_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_l8 : unsigned(7 downto 0);
variable REG_VAR_current_deo_phase : unsigned(7 downto 0);
variable REG_VAR_deo_param0 : unsigned(7 downto 0);
variable REG_VAR_deo_param1 : unsigned(7 downto 0);
variable REG_VAR_is_second_deo : unsigned(0 downto 0);
variable REG_VAR_is_phase_3 : unsigned(0 downto 0);
variable REG_VAR_is_phase_4 : unsigned(0 downto 0);
variable REG_VAR_result : opcode_result_t;
variable REG_VAR_device_out_result : device_out_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_l8 := l8;
  REG_VAR_current_deo_phase := current_deo_phase;
  REG_VAR_deo_param0 := deo_param0;
  REG_VAR_deo_param1 := deo_param1;
  REG_VAR_is_second_deo := is_second_deo;
  REG_VAR_is_phase_3 := is_phase_3;
  REG_VAR_is_phase_4 := is_phase_4;
  REG_VAR_result := result;
  REG_VAR_device_out_result := device_out_result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_current_deo_phase_uxn_opcodes_h_l546_c3_3298 := resize(to_unsigned(0, 1), 8);
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_iftrue := VAR_current_deo_phase_uxn_opcodes_h_l546_c3_3298;
     VAR_sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l549_c3_9a1e := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l549_c3_9a1e;
     VAR_MUX_uxn_opcodes_h_l557_c17_bfc8_iffalse := to_unsigned(0, 1);
     VAR_is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_iftrue := to_unsigned(0, 1);
     VAR_current_deo_phase_uxn_opcodes_h_l572_c4_b061 := resize(to_unsigned(0, 1), 8);
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_iftrue := VAR_current_deo_phase_uxn_opcodes_h_l572_c4_b061;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_right := to_unsigned(0, 1);
     VAR_is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l552_c3_f51c := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l552_c3_f51c;
     VAR_MUX_uxn_opcodes_h_l557_c17_bfc8_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l557_c17_c8c7_right := to_unsigned(4, 3);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l543_c3_51f3 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l543_c3_51f3;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_iftrue := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l556_c17_aaf6_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_y := resize(to_signed(-3, 3), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_right := to_unsigned(2, 2);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l560_c32_60a0_right := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l556_c17_aaf6_iffalse := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l562_c30_d095_iffalse := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c17_5fcc_right := to_unsigned(3, 2);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l575_c4_0ea3_right := to_unsigned(1, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_device_ram_read := previous_device_ram_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l575_c4_0ea3_left := current_deo_phase;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue := current_deo_phase;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_iftrue := current_deo_phase;
     VAR_device_out_uxn_opcodes_h_l563_c23_d468_phase := current_deo_phase;
     VAR_deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_iftrue := deo_param0;
     VAR_deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue := deo_param0;
     VAR_deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_iftrue := deo_param0;
     VAR_deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_iftrue := deo_param1;
     VAR_deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue := deo_param1;
     VAR_deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_iftrue := deo_param1;
     VAR_device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_iftrue := device_out_result;
     VAR_device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue := device_out_result;
     VAR_device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_iftrue := device_out_result;
     VAR_sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_ins := VAR_ins;
     VAR_is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_iftrue := is_phase_3;
     VAR_is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue := is_phase_3;
     VAR_is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_iftrue := is_phase_3;
     VAR_is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_iftrue := is_phase_4;
     VAR_is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue := is_phase_4;
     VAR_is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_iftrue := is_phase_4;
     VAR_BIN_OP_AND_uxn_opcodes_h_l570_c24_c405_right := is_second_deo;
     VAR_MUX_uxn_opcodes_h_l560_c16_ee8b_cond := is_second_deo;
     VAR_MUX_uxn_opcodes_h_l561_c16_e93e_cond := is_second_deo;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue := is_second_deo;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_iftrue := is_second_deo;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_iffalse := is_second_deo;
     VAR_MUX_uxn_opcodes_h_l558_c8_9c1c_iffalse := l8;
     VAR_l8_MUX_uxn_opcodes_h_l539_c2_8124_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l551_c7_205d_iftrue := l8;
     VAR_MUX_uxn_opcodes_h_l559_c8_9d6a_iffalse := n8;
     VAR_n8_MUX_uxn_opcodes_h_l539_c2_8124_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l551_c7_205d_iftrue := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c17_5fcc_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l557_c17_c8c7_left := VAR_phase;
     VAR_device_out_uxn_opcodes_h_l563_c23_d468_previous_device_ram_read := VAR_previous_device_ram_read;
     VAR_device_out_uxn_opcodes_h_l563_c23_d468_previous_ram_read := VAR_previous_ram_read;
     VAR_MUX_uxn_opcodes_h_l558_c8_9c1c_iftrue := VAR_previous_stack_read;
     VAR_MUX_uxn_opcodes_h_l559_c8_9d6a_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l551_c7_205d_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l560_c32_60a0_left := t8;
     VAR_MUX_uxn_opcodes_h_l560_c16_ee8b_iffalse := t8;
     VAR_t8_MUX_uxn_opcodes_h_l539_c2_8124_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l551_c7_205d_iffalse := t8;
     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_85a2 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_85a2_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_127b LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_127b_return_output := result.u16_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_271a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_271a_return_output := result.is_device_ram_write;

     -- sp_relative_shift[uxn_opcodes_h_l562_c43_1dbf] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_ins;
     sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_x <= VAR_sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_x;
     sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_y <= VAR_sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_return_output := sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l557_c17_c8c7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l557_c17_c8c7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l557_c17_c8c7_left;
     BIN_OP_EQ_uxn_opcodes_h_l557_c17_c8c7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l557_c17_c8c7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l557_c17_c8c7_return_output := BIN_OP_EQ_uxn_opcodes_h_l557_c17_c8c7_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l551_c7_205d] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l551_c7_205d_return_output := result.stack_address_sp_offset;

     -- BIN_OP_PLUS[uxn_opcodes_h_l560_c32_60a0] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l560_c32_60a0_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l560_c32_60a0_left;
     BIN_OP_PLUS_uxn_opcodes_h_l560_c32_60a0_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l560_c32_60a0_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l560_c32_60a0_return_output := BIN_OP_PLUS_uxn_opcodes_h_l560_c32_60a0_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_4e2e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_4e2e_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_c949 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_c949_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l548_c11_6174] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_left;
     BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output := BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l539_c6_9f48] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_left;
     BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output := BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_8fa6 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_8fa6_return_output := result.device_ram_address;

     -- BIN_OP_EQ[uxn_opcodes_h_l551_c11_ffc2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_left;
     BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output := BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l556_c17_5fcc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l556_c17_5fcc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c17_5fcc_left;
     BIN_OP_EQ_uxn_opcodes_h_l556_c17_5fcc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c17_5fcc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c17_5fcc_return_output := BIN_OP_EQ_uxn_opcodes_h_l556_c17_5fcc_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l548_l551_DUPLICATE_336e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l548_l551_DUPLICATE_336e_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_176c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_176c_return_output := result.vram_write_layer;

     -- BIN_OP_PLUS[uxn_opcodes_h_l575_c4_0ea3] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l575_c4_0ea3_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l575_c4_0ea3_left;
     BIN_OP_PLUS_uxn_opcodes_h_l575_c4_0ea3_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l575_c4_0ea3_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l575_c4_0ea3_return_output := BIN_OP_PLUS_uxn_opcodes_h_l575_c4_0ea3_return_output;

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output;
     VAR_deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output;
     VAR_deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output;
     VAR_is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output;
     VAR_is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l539_c2_8124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l539_c2_8124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l539_c2_8124_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l539_c6_9f48_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output;
     VAR_deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output;
     VAR_deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output;
     VAR_is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output;
     VAR_is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l548_c7_ce40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l548_c7_ce40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l548_c7_ce40_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l548_c11_6174_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output;
     VAR_deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output;
     VAR_deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output;
     VAR_is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output;
     VAR_is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l551_c7_205d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l551_c7_205d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l551_c7_205d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l551_c11_ffc2_return_output;
     VAR_MUX_uxn_opcodes_h_l556_c17_aaf6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l556_c17_5fcc_return_output;
     VAR_MUX_uxn_opcodes_h_l557_c17_bfc8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l557_c17_c8c7_return_output;
     VAR_MUX_uxn_opcodes_h_l560_c16_ee8b_iftrue := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l560_c32_60a0_return_output, 8);
     VAR_current_deo_phase_uxn_opcodes_h_l575_c4_f6a7 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l575_c4_0ea3_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_85a2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_85a2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_85a2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_127b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_127b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_127b_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_271a_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_271a_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_271a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l548_l551_DUPLICATE_336e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l548_l551_DUPLICATE_336e_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_c949_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_c949_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_c949_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_176c_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_176c_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_176c_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_8fa6_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_8fa6_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_8fa6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_4e2e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_4e2e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l548_l551_l539_DUPLICATE_4e2e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l551_c7_205d_return_output;
     VAR_MUX_uxn_opcodes_h_l562_c30_d095_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l562_c43_1dbf_return_output;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_iffalse := VAR_current_deo_phase_uxn_opcodes_h_l575_c4_f6a7;
     -- MUX[uxn_opcodes_h_l556_c17_aaf6] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l556_c17_aaf6_cond <= VAR_MUX_uxn_opcodes_h_l556_c17_aaf6_cond;
     MUX_uxn_opcodes_h_l556_c17_aaf6_iftrue <= VAR_MUX_uxn_opcodes_h_l556_c17_aaf6_iftrue;
     MUX_uxn_opcodes_h_l556_c17_aaf6_iffalse <= VAR_MUX_uxn_opcodes_h_l556_c17_aaf6_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l556_c17_aaf6_return_output := MUX_uxn_opcodes_h_l556_c17_aaf6_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l548_c7_ce40] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l551_c7_205d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_return_output;

     -- t8_MUX[uxn_opcodes_h_l551_c7_205d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l551_c7_205d_cond <= VAR_t8_MUX_uxn_opcodes_h_l551_c7_205d_cond;
     t8_MUX_uxn_opcodes_h_l551_c7_205d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l551_c7_205d_iftrue;
     t8_MUX_uxn_opcodes_h_l551_c7_205d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l551_c7_205d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l551_c7_205d_return_output := t8_MUX_uxn_opcodes_h_l551_c7_205d_return_output;

     -- MUX[uxn_opcodes_h_l560_c16_ee8b] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l560_c16_ee8b_cond <= VAR_MUX_uxn_opcodes_h_l560_c16_ee8b_cond;
     MUX_uxn_opcodes_h_l560_c16_ee8b_iftrue <= VAR_MUX_uxn_opcodes_h_l560_c16_ee8b_iftrue;
     MUX_uxn_opcodes_h_l560_c16_ee8b_iffalse <= VAR_MUX_uxn_opcodes_h_l560_c16_ee8b_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l560_c16_ee8b_return_output := MUX_uxn_opcodes_h_l560_c16_ee8b_return_output;

     -- MUX[uxn_opcodes_h_l557_c17_bfc8] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l557_c17_bfc8_cond <= VAR_MUX_uxn_opcodes_h_l557_c17_bfc8_cond;
     MUX_uxn_opcodes_h_l557_c17_bfc8_iftrue <= VAR_MUX_uxn_opcodes_h_l557_c17_bfc8_iftrue;
     MUX_uxn_opcodes_h_l557_c17_bfc8_iffalse <= VAR_MUX_uxn_opcodes_h_l557_c17_bfc8_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l557_c17_bfc8_return_output := MUX_uxn_opcodes_h_l557_c17_bfc8_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;
     VAR_MUX_uxn_opcodes_h_l558_c8_9c1c_cond := VAR_MUX_uxn_opcodes_h_l556_c17_aaf6_return_output;
     VAR_MUX_uxn_opcodes_h_l562_c30_d095_cond := VAR_MUX_uxn_opcodes_h_l556_c17_aaf6_return_output;
     VAR_is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_iffalse := VAR_MUX_uxn_opcodes_h_l556_c17_aaf6_return_output;
     VAR_MUX_uxn_opcodes_h_l559_c8_9d6a_cond := VAR_MUX_uxn_opcodes_h_l557_c17_bfc8_return_output;
     VAR_is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_iffalse := VAR_MUX_uxn_opcodes_h_l557_c17_bfc8_return_output;
     VAR_deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_iffalse := VAR_MUX_uxn_opcodes_h_l560_c16_ee8b_return_output;
     VAR_device_out_uxn_opcodes_h_l563_c23_d468_device_address := VAR_MUX_uxn_opcodes_h_l560_c16_ee8b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l551_c7_205d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse := VAR_t8_MUX_uxn_opcodes_h_l551_c7_205d_return_output;
     -- t8_MUX[uxn_opcodes_h_l548_c7_ce40] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l548_c7_ce40_cond <= VAR_t8_MUX_uxn_opcodes_h_l548_c7_ce40_cond;
     t8_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue;
     t8_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l548_c7_ce40_return_output := t8_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;

     -- MUX[uxn_opcodes_h_l559_c8_9d6a] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l559_c8_9d6a_cond <= VAR_MUX_uxn_opcodes_h_l559_c8_9d6a_cond;
     MUX_uxn_opcodes_h_l559_c8_9d6a_iftrue <= VAR_MUX_uxn_opcodes_h_l559_c8_9d6a_iftrue;
     MUX_uxn_opcodes_h_l559_c8_9d6a_iffalse <= VAR_MUX_uxn_opcodes_h_l559_c8_9d6a_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l559_c8_9d6a_return_output := MUX_uxn_opcodes_h_l559_c8_9d6a_return_output;

     -- MUX[uxn_opcodes_h_l562_c30_d095] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l562_c30_d095_cond <= VAR_MUX_uxn_opcodes_h_l562_c30_d095_cond;
     MUX_uxn_opcodes_h_l562_c30_d095_iftrue <= VAR_MUX_uxn_opcodes_h_l562_c30_d095_iftrue;
     MUX_uxn_opcodes_h_l562_c30_d095_iffalse <= VAR_MUX_uxn_opcodes_h_l562_c30_d095_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l562_c30_d095_return_output := MUX_uxn_opcodes_h_l562_c30_d095_return_output;

     -- is_phase_4_MUX[uxn_opcodes_h_l551_c7_205d] LATENCY=0
     -- Inputs
     is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_cond <= VAR_is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_cond;
     is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_iftrue <= VAR_is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_iftrue;
     is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_iffalse <= VAR_is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_iffalse;
     -- Outputs
     VAR_is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_return_output := is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_return_output;

     -- deo_param0_MUX[uxn_opcodes_h_l551_c7_205d] LATENCY=0
     -- Inputs
     deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_cond <= VAR_deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_cond;
     deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_iftrue <= VAR_deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_iftrue;
     deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_iffalse <= VAR_deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_iffalse;
     -- Outputs
     VAR_deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_return_output := deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_return_output;

     -- is_phase_3_MUX[uxn_opcodes_h_l551_c7_205d] LATENCY=0
     -- Inputs
     is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_cond <= VAR_is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_cond;
     is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_iftrue <= VAR_is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_iftrue;
     is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_iffalse <= VAR_is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_iffalse;
     -- Outputs
     VAR_is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_return_output := is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_return_output;

     -- MUX[uxn_opcodes_h_l558_c8_9c1c] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l558_c8_9c1c_cond <= VAR_MUX_uxn_opcodes_h_l558_c8_9c1c_cond;
     MUX_uxn_opcodes_h_l558_c8_9c1c_iftrue <= VAR_MUX_uxn_opcodes_h_l558_c8_9c1c_iftrue;
     MUX_uxn_opcodes_h_l558_c8_9c1c_iffalse <= VAR_MUX_uxn_opcodes_h_l558_c8_9c1c_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l558_c8_9c1c_return_output := MUX_uxn_opcodes_h_l558_c8_9c1c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l548_c7_ce40] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l551_c7_205d] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_return_output;

     -- Submodule level 3
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l551_c7_205d_return_output;
     VAR_MUX_uxn_opcodes_h_l561_c16_e93e_iffalse := VAR_MUX_uxn_opcodes_h_l558_c8_9c1c_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l551_c7_205d_iffalse := VAR_MUX_uxn_opcodes_h_l558_c8_9c1c_return_output;
     VAR_MUX_uxn_opcodes_h_l561_c16_e93e_iftrue := VAR_MUX_uxn_opcodes_h_l559_c8_9d6a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l551_c7_205d_iffalse := VAR_MUX_uxn_opcodes_h_l559_c8_9d6a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_iffalse := VAR_MUX_uxn_opcodes_h_l562_c30_d095_return_output;
     VAR_deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse := VAR_deo_param0_MUX_uxn_opcodes_h_l551_c7_205d_return_output;
     VAR_is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse := VAR_is_phase_3_MUX_uxn_opcodes_h_l551_c7_205d_return_output;
     VAR_is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse := VAR_is_phase_4_MUX_uxn_opcodes_h_l551_c7_205d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l539_c2_8124_iffalse := VAR_t8_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;
     -- n8_MUX[uxn_opcodes_h_l551_c7_205d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l551_c7_205d_cond <= VAR_n8_MUX_uxn_opcodes_h_l551_c7_205d_cond;
     n8_MUX_uxn_opcodes_h_l551_c7_205d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l551_c7_205d_iftrue;
     n8_MUX_uxn_opcodes_h_l551_c7_205d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l551_c7_205d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l551_c7_205d_return_output := n8_MUX_uxn_opcodes_h_l551_c7_205d_return_output;

     -- is_phase_3_MUX[uxn_opcodes_h_l548_c7_ce40] LATENCY=0
     -- Inputs
     is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_cond <= VAR_is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_cond;
     is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue <= VAR_is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue;
     is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse <= VAR_is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse;
     -- Outputs
     VAR_is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_return_output := is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;

     -- l8_MUX[uxn_opcodes_h_l551_c7_205d] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l551_c7_205d_cond <= VAR_l8_MUX_uxn_opcodes_h_l551_c7_205d_cond;
     l8_MUX_uxn_opcodes_h_l551_c7_205d_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l551_c7_205d_iftrue;
     l8_MUX_uxn_opcodes_h_l551_c7_205d_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l551_c7_205d_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l551_c7_205d_return_output := l8_MUX_uxn_opcodes_h_l551_c7_205d_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l555_c1_b0c5] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l551_c7_205d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_return_output;

     -- deo_param0_MUX[uxn_opcodes_h_l548_c7_ce40] LATENCY=0
     -- Inputs
     deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_cond <= VAR_deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_cond;
     deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue <= VAR_deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue;
     deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse <= VAR_deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse;
     -- Outputs
     VAR_deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_return_output := deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;

     -- t8_MUX[uxn_opcodes_h_l539_c2_8124] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l539_c2_8124_cond <= VAR_t8_MUX_uxn_opcodes_h_l539_c2_8124_cond;
     t8_MUX_uxn_opcodes_h_l539_c2_8124_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l539_c2_8124_iftrue;
     t8_MUX_uxn_opcodes_h_l539_c2_8124_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l539_c2_8124_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l539_c2_8124_return_output := t8_MUX_uxn_opcodes_h_l539_c2_8124_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l539_c2_8124] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_return_output;

     -- is_phase_4_MUX[uxn_opcodes_h_l548_c7_ce40] LATENCY=0
     -- Inputs
     is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_cond <= VAR_is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_cond;
     is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue <= VAR_is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue;
     is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse <= VAR_is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse;
     -- Outputs
     VAR_is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_return_output := is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;

     -- MUX[uxn_opcodes_h_l561_c16_e93e] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l561_c16_e93e_cond <= VAR_MUX_uxn_opcodes_h_l561_c16_e93e_cond;
     MUX_uxn_opcodes_h_l561_c16_e93e_iftrue <= VAR_MUX_uxn_opcodes_h_l561_c16_e93e_iftrue;
     MUX_uxn_opcodes_h_l561_c16_e93e_iffalse <= VAR_MUX_uxn_opcodes_h_l561_c16_e93e_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l561_c16_e93e_return_output := MUX_uxn_opcodes_h_l561_c16_e93e_return_output;

     -- Submodule level 4
     VAR_device_out_uxn_opcodes_h_l563_c23_d468_CLOCK_ENABLE := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l555_c1_b0c5_return_output;
     VAR_deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_iffalse := VAR_MUX_uxn_opcodes_h_l561_c16_e93e_return_output;
     VAR_device_out_uxn_opcodes_h_l563_c23_d468_value := VAR_MUX_uxn_opcodes_h_l561_c16_e93e_return_output;
     VAR_deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_iffalse := VAR_deo_param0_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;
     VAR_is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_iffalse := VAR_is_phase_3_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;
     VAR_is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_iffalse := VAR_is_phase_4_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse := VAR_l8_MUX_uxn_opcodes_h_l551_c7_205d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse := VAR_n8_MUX_uxn_opcodes_h_l551_c7_205d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l551_c7_205d_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l539_c2_8124_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l548_c7_ce40] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;

     -- is_phase_3_MUX[uxn_opcodes_h_l539_c2_8124] LATENCY=0
     -- Inputs
     is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_cond <= VAR_is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_cond;
     is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_iftrue <= VAR_is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_iftrue;
     is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_iffalse <= VAR_is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_iffalse;
     -- Outputs
     VAR_is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_return_output := is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_return_output;

     -- device_out[uxn_opcodes_h_l563_c23_d468] LATENCY=0
     -- Clock enable
     device_out_uxn_opcodes_h_l563_c23_d468_CLOCK_ENABLE <= VAR_device_out_uxn_opcodes_h_l563_c23_d468_CLOCK_ENABLE;
     -- Inputs
     device_out_uxn_opcodes_h_l563_c23_d468_device_address <= VAR_device_out_uxn_opcodes_h_l563_c23_d468_device_address;
     device_out_uxn_opcodes_h_l563_c23_d468_value <= VAR_device_out_uxn_opcodes_h_l563_c23_d468_value;
     device_out_uxn_opcodes_h_l563_c23_d468_phase <= VAR_device_out_uxn_opcodes_h_l563_c23_d468_phase;
     device_out_uxn_opcodes_h_l563_c23_d468_previous_device_ram_read <= VAR_device_out_uxn_opcodes_h_l563_c23_d468_previous_device_ram_read;
     device_out_uxn_opcodes_h_l563_c23_d468_previous_ram_read <= VAR_device_out_uxn_opcodes_h_l563_c23_d468_previous_ram_read;
     -- Outputs
     VAR_device_out_uxn_opcodes_h_l563_c23_d468_return_output := device_out_uxn_opcodes_h_l563_c23_d468_return_output;

     -- is_phase_4_MUX[uxn_opcodes_h_l539_c2_8124] LATENCY=0
     -- Inputs
     is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_cond <= VAR_is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_cond;
     is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_iftrue <= VAR_is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_iftrue;
     is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_iffalse <= VAR_is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_iffalse;
     -- Outputs
     VAR_is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_return_output := is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_return_output;

     -- l8_MUX[uxn_opcodes_h_l548_c7_ce40] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l548_c7_ce40_cond <= VAR_l8_MUX_uxn_opcodes_h_l548_c7_ce40_cond;
     l8_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue;
     l8_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l548_c7_ce40_return_output := l8_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;

     -- deo_param0_MUX[uxn_opcodes_h_l539_c2_8124] LATENCY=0
     -- Inputs
     deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_cond <= VAR_deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_cond;
     deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_iftrue <= VAR_deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_iftrue;
     deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_iffalse <= VAR_deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_iffalse;
     -- Outputs
     VAR_deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_return_output := deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_return_output;

     -- deo_param1_MUX[uxn_opcodes_h_l551_c7_205d] LATENCY=0
     -- Inputs
     deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_cond <= VAR_deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_cond;
     deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_iftrue <= VAR_deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_iftrue;
     deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_iffalse <= VAR_deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_iffalse;
     -- Outputs
     VAR_deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_return_output := deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_return_output;

     -- n8_MUX[uxn_opcodes_h_l548_c7_ce40] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l548_c7_ce40_cond <= VAR_n8_MUX_uxn_opcodes_h_l548_c7_ce40_cond;
     n8_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue;
     n8_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l548_c7_ce40_return_output := n8_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;

     -- Submodule level 5
     REG_VAR_deo_param0 := VAR_deo_param0_MUX_uxn_opcodes_h_l539_c2_8124_return_output;
     VAR_deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse := VAR_deo_param1_MUX_uxn_opcodes_h_l551_c7_205d_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_iffalse := VAR_device_out_uxn_opcodes_h_l563_c23_d468_return_output;
     REG_VAR_is_phase_3 := VAR_is_phase_3_MUX_uxn_opcodes_h_l539_c2_8124_return_output;
     REG_VAR_is_phase_4 := VAR_is_phase_4_MUX_uxn_opcodes_h_l539_c2_8124_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l539_c2_8124_iffalse := VAR_l8_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l539_c2_8124_iffalse := VAR_n8_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;
     -- CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d_uxn_opcodes_h_l570_l571_DUPLICATE_f81b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d_uxn_opcodes_h_l570_l571_DUPLICATE_f81b_return_output := VAR_device_out_uxn_opcodes_h_l563_c23_d468_return_output.is_deo_done;

     -- device_out_result_MUX[uxn_opcodes_h_l551_c7_205d] LATENCY=0
     -- Inputs
     device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_cond <= VAR_device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_cond;
     device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_iftrue <= VAR_device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_iftrue;
     device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_iffalse <= VAR_device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_iffalse;
     -- Outputs
     VAR_device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_return_output := device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_return_output;

     -- CONST_REF_RD_uint1_t_device_out_result_t_is_vram_write_d41d[uxn_opcodes_h_l566_c26_75a1] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_vram_write_d41d_uxn_opcodes_h_l566_c26_75a1_return_output := VAR_device_out_uxn_opcodes_h_l563_c23_d468_return_output.is_vram_write;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l539_c2_8124] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_return_output;

     -- l8_MUX[uxn_opcodes_h_l539_c2_8124] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l539_c2_8124_cond <= VAR_l8_MUX_uxn_opcodes_h_l539_c2_8124_cond;
     l8_MUX_uxn_opcodes_h_l539_c2_8124_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l539_c2_8124_iftrue;
     l8_MUX_uxn_opcodes_h_l539_c2_8124_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l539_c2_8124_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l539_c2_8124_return_output := l8_MUX_uxn_opcodes_h_l539_c2_8124_return_output;

     -- n8_MUX[uxn_opcodes_h_l539_c2_8124] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l539_c2_8124_cond <= VAR_n8_MUX_uxn_opcodes_h_l539_c2_8124_cond;
     n8_MUX_uxn_opcodes_h_l539_c2_8124_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l539_c2_8124_iftrue;
     n8_MUX_uxn_opcodes_h_l539_c2_8124_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l539_c2_8124_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l539_c2_8124_return_output := n8_MUX_uxn_opcodes_h_l539_c2_8124_return_output;

     -- CONST_REF_RD_uint1_t_device_out_result_t_vram_write_layer_d41d[uxn_opcodes_h_l567_c29_f9a5] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_out_result_t_vram_write_layer_d41d_uxn_opcodes_h_l567_c29_f9a5_return_output := VAR_device_out_uxn_opcodes_h_l563_c23_d468_return_output.vram_write_layer;

     -- CONST_REF_RD_uint8_t_device_out_result_t_u8_value_d41d[uxn_opcodes_h_l569_c21_f77c] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_out_result_t_u8_value_d41d_uxn_opcodes_h_l569_c21_f77c_return_output := VAR_device_out_uxn_opcodes_h_l563_c23_d468_return_output.u8_value;

     -- CONST_REF_RD_uint1_t_device_out_result_t_is_device_ram_write_d41d[uxn_opcodes_h_l564_c32_f2a0] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l564_c32_f2a0_return_output := VAR_device_out_uxn_opcodes_h_l563_c23_d468_return_output.is_device_ram_write;

     -- CONST_REF_RD_uint8_t_device_out_result_t_device_ram_address_d41d[uxn_opcodes_h_l565_c31_6b03] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_out_result_t_device_ram_address_d41d_uxn_opcodes_h_l565_c31_6b03_return_output := VAR_device_out_uxn_opcodes_h_l563_c23_d468_return_output.device_ram_address;

     -- CONST_REF_RD_uint16_t_device_out_result_t_u16_addr_d41d[uxn_opcodes_h_l568_c22_b6cb] LATENCY=0
     VAR_CONST_REF_RD_uint16_t_device_out_result_t_u16_addr_d41d_uxn_opcodes_h_l568_c22_b6cb_return_output := VAR_device_out_uxn_opcodes_h_l563_c23_d468_return_output.u16_addr;

     -- deo_param1_MUX[uxn_opcodes_h_l548_c7_ce40] LATENCY=0
     -- Inputs
     deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_cond <= VAR_deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_cond;
     deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue <= VAR_deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue;
     deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse <= VAR_deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse;
     -- Outputs
     VAR_deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_return_output := deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;

     -- Submodule level 6
     VAR_result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_iffalse := VAR_CONST_REF_RD_uint16_t_device_out_result_t_u16_addr_d41d_uxn_opcodes_h_l568_c22_b6cb_return_output;
     VAR_BIN_OP_AND_uxn_opcodes_h_l570_c24_c405_left := VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d_uxn_opcodes_h_l570_l571_DUPLICATE_f81b_return_output;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_cond := VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d_uxn_opcodes_h_l570_l571_DUPLICATE_f81b_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_cond := VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d_uxn_opcodes_h_l570_l571_DUPLICATE_f81b_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_iffalse := VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l564_c32_f2a0_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_iffalse := VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_vram_write_d41d_uxn_opcodes_h_l566_c26_75a1_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_iffalse := VAR_CONST_REF_RD_uint1_t_device_out_result_t_vram_write_layer_d41d_uxn_opcodes_h_l567_c29_f9a5_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_iffalse := VAR_CONST_REF_RD_uint8_t_device_out_result_t_device_ram_address_d41d_uxn_opcodes_h_l565_c31_6b03_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_iffalse := VAR_CONST_REF_RD_uint8_t_device_out_result_t_u8_value_d41d_uxn_opcodes_h_l569_c21_f77c_return_output;
     VAR_deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_iffalse := VAR_deo_param1_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse := VAR_device_out_result_MUX_uxn_opcodes_h_l551_c7_205d_return_output;
     REG_VAR_l8 := VAR_l8_MUX_uxn_opcodes_h_l539_c2_8124_return_output;
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l539_c2_8124_return_output;
     -- result_device_ram_address_MUX[uxn_opcodes_h_l551_c7_205d] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_return_output;

     -- current_deo_phase_MUX[uxn_opcodes_h_l571_c3_6837] LATENCY=0
     -- Inputs
     current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_cond <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_cond;
     current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_iftrue <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_iftrue;
     current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_iffalse <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_iffalse;
     -- Outputs
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_return_output := current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l551_c7_205d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_return_output := result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l551_c7_205d] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l551_c7_205d] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_cond;
     result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_return_output := result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_return_output;

     -- deo_param1_MUX[uxn_opcodes_h_l539_c2_8124] LATENCY=0
     -- Inputs
     deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_cond <= VAR_deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_cond;
     deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_iftrue <= VAR_deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_iftrue;
     deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_iffalse <= VAR_deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_iffalse;
     -- Outputs
     VAR_deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_return_output := deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_return_output;

     -- result_vram_write_layer_MUX[uxn_opcodes_h_l551_c7_205d] LATENCY=0
     -- Inputs
     result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_cond <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_cond;
     result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_iftrue <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_iftrue;
     result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_iffalse <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_iffalse;
     -- Outputs
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_return_output := result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l570_c24_c405] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l570_c24_c405_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l570_c24_c405_left;
     BIN_OP_AND_uxn_opcodes_h_l570_c24_c405_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l570_c24_c405_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l570_c24_c405_return_output := BIN_OP_AND_uxn_opcodes_h_l570_c24_c405_return_output;

     -- device_out_result_MUX[uxn_opcodes_h_l548_c7_ce40] LATENCY=0
     -- Inputs
     device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_cond <= VAR_device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_cond;
     device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue <= VAR_device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue;
     device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse <= VAR_device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse;
     -- Outputs
     VAR_device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_return_output := device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;

     -- result_is_device_ram_write_MUX[uxn_opcodes_h_l551_c7_205d] LATENCY=0
     -- Inputs
     result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_cond <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_cond;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_iftrue <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_iftrue;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_iffalse <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_iffalse;
     -- Outputs
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_return_output := result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_return_output;

     -- is_second_deo_MUX[uxn_opcodes_h_l571_c3_6837] LATENCY=0
     -- Inputs
     is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_cond <= VAR_is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_cond;
     is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_iftrue <= VAR_is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_iftrue;
     is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_iffalse <= VAR_is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_iffalse;
     -- Outputs
     VAR_is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_return_output := is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_return_output;

     -- Submodule level 7
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_iffalse := VAR_BIN_OP_AND_uxn_opcodes_h_l570_c24_c405_return_output;
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_iffalse := VAR_current_deo_phase_MUX_uxn_opcodes_h_l571_c3_6837_return_output;
     REG_VAR_deo_param1 := VAR_deo_param1_MUX_uxn_opcodes_h_l539_c2_8124_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_iffalse := VAR_device_out_result_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_iffalse := VAR_is_second_deo_MUX_uxn_opcodes_h_l571_c3_6837_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l551_c7_205d_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse := VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l551_c7_205d_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse := VAR_result_is_vram_write_MUX_uxn_opcodes_h_l551_c7_205d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l551_c7_205d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l551_c7_205d_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse := VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l551_c7_205d_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l551_c7_205d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l548_c7_ce40] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_cond;
     result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_return_output := result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;

     -- result_vram_write_layer_MUX[uxn_opcodes_h_l548_c7_ce40] LATENCY=0
     -- Inputs
     result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_cond <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_cond;
     result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue;
     result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse;
     -- Outputs
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_return_output := result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l548_c7_ce40] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_cond;
     result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_return_output := result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;

     -- current_deo_phase_MUX[uxn_opcodes_h_l551_c7_205d] LATENCY=0
     -- Inputs
     current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_cond <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_cond;
     current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_iftrue <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_iftrue;
     current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_iffalse <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_iffalse;
     -- Outputs
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_return_output := current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_return_output;

     -- is_second_deo_MUX[uxn_opcodes_h_l551_c7_205d] LATENCY=0
     -- Inputs
     is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_cond <= VAR_is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_cond;
     is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_iftrue <= VAR_is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_iftrue;
     is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_iffalse <= VAR_is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_iffalse;
     -- Outputs
     VAR_is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_return_output := is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l548_c7_ce40] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;

     -- result_is_device_ram_write_MUX[uxn_opcodes_h_l548_c7_ce40] LATENCY=0
     -- Inputs
     result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_cond <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_cond;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse;
     -- Outputs
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_return_output := result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;

     -- device_out_result_MUX[uxn_opcodes_h_l539_c2_8124] LATENCY=0
     -- Inputs
     device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_cond <= VAR_device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_cond;
     device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_iftrue <= VAR_device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_iftrue;
     device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_iffalse <= VAR_device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_iffalse;
     -- Outputs
     VAR_device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_return_output := device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_return_output;

     -- result_device_ram_address_MUX[uxn_opcodes_h_l548_c7_ce40] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;

     -- Submodule level 8
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse := VAR_current_deo_phase_MUX_uxn_opcodes_h_l551_c7_205d_return_output;
     REG_VAR_device_out_result := VAR_device_out_result_MUX_uxn_opcodes_h_l539_c2_8124_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse := VAR_is_second_deo_MUX_uxn_opcodes_h_l551_c7_205d_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_iffalse := VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l551_c7_205d_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_iffalse := VAR_result_is_vram_write_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_iffalse := VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l548_c7_ce40] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l539_c2_8124] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_cond;
     result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_return_output := result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_return_output;

     -- result_device_ram_address_MUX[uxn_opcodes_h_l539_c2_8124] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_return_output;

     -- current_deo_phase_MUX[uxn_opcodes_h_l548_c7_ce40] LATENCY=0
     -- Inputs
     current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_cond <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_cond;
     current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue;
     current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse;
     -- Outputs
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_return_output := current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;

     -- result_vram_write_layer_MUX[uxn_opcodes_h_l539_c2_8124] LATENCY=0
     -- Inputs
     result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_cond <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_cond;
     result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_iftrue <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_iftrue;
     result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_iffalse <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_iffalse;
     -- Outputs
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_return_output := result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_return_output;

     -- result_is_device_ram_write_MUX[uxn_opcodes_h_l539_c2_8124] LATENCY=0
     -- Inputs
     result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_cond <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_cond;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_iftrue <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_iftrue;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_iffalse <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_iffalse;
     -- Outputs
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_return_output := result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l539_c2_8124] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_cond;
     result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_return_output := result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_return_output;

     -- is_second_deo_MUX[uxn_opcodes_h_l548_c7_ce40] LATENCY=0
     -- Inputs
     is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_cond <= VAR_is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_cond;
     is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue <= VAR_is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_iftrue;
     is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse <= VAR_is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_iffalse;
     -- Outputs
     VAR_is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_return_output := is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l539_c2_8124] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_return_output;

     -- Submodule level 9
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_iffalse := VAR_current_deo_phase_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;
     VAR_is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_iffalse := VAR_is_second_deo_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l548_c7_ce40_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l539_c2_8124] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_return_output;

     -- is_second_deo_MUX[uxn_opcodes_h_l539_c2_8124] LATENCY=0
     -- Inputs
     is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_cond <= VAR_is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_cond;
     is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_iftrue <= VAR_is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_iftrue;
     is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_iffalse <= VAR_is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_iffalse;
     -- Outputs
     VAR_is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_return_output := is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_return_output;

     -- current_deo_phase_MUX[uxn_opcodes_h_l539_c2_8124] LATENCY=0
     -- Inputs
     current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_cond <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_cond;
     current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_iftrue <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_iftrue;
     current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_iffalse <= VAR_current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_iffalse;
     -- Outputs
     VAR_current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_return_output := current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_return_output;

     -- Submodule level 10
     REG_VAR_current_deo_phase := VAR_current_deo_phase_MUX_uxn_opcodes_h_l539_c2_8124_return_output;
     REG_VAR_is_second_deo := VAR_is_second_deo_MUX_uxn_opcodes_h_l539_c2_8124_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_f18e_uxn_opcodes_h_l579_l533_DUPLICATE_d422 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_f18e_uxn_opcodes_h_l579_l533_DUPLICATE_d422_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_f18e(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l539_c2_8124_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l539_c2_8124_return_output);

     -- Submodule level 11
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_f18e_uxn_opcodes_h_l579_l533_DUPLICATE_d422_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_f18e_uxn_opcodes_h_l579_l533_DUPLICATE_d422_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_l8 <= REG_VAR_l8;
REG_COMB_current_deo_phase <= REG_VAR_current_deo_phase;
REG_COMB_deo_param0 <= REG_VAR_deo_param0;
REG_COMB_deo_param1 <= REG_VAR_deo_param1;
REG_COMB_is_second_deo <= REG_VAR_is_second_deo;
REG_COMB_is_phase_3 <= REG_VAR_is_phase_3;
REG_COMB_is_phase_4 <= REG_VAR_is_phase_4;
REG_COMB_result <= REG_VAR_result;
REG_COMB_device_out_result <= REG_VAR_device_out_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     l8 <= REG_COMB_l8;
     current_deo_phase <= REG_COMB_current_deo_phase;
     deo_param0 <= REG_COMB_deo_param0;
     deo_param1 <= REG_COMB_deo_param1;
     is_second_deo <= REG_COMB_is_second_deo;
     is_phase_3 <= REG_COMB_is_phase_3;
     is_phase_4 <= REG_COMB_is_phase_4;
     result <= REG_COMB_result;
     device_out_result <= REG_COMB_device_out_result;
 end if;
 end if;
end process;

end arch;
