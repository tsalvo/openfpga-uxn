-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity gth_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end gth_0CLK_226c8821;
architecture arch of gth_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1832_c6_9abb]
signal BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1832_c2_0399]
signal t8_MUX_uxn_opcodes_h_l1832_c2_0399_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1832_c2_0399_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1832_c2_0399]
signal n8_MUX_uxn_opcodes_h_l1832_c2_0399_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1832_c2_0399_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1832_c2_0399]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1832_c2_0399]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1832_c2_0399]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1832_c2_0399]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1832_c2_0399]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1832_c2_0399]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1832_c2_0399]
signal result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1832_c2_0399]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1832_c2_0399]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1845_c11_726c]
signal BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1845_c7_9f69]
signal t8_MUX_uxn_opcodes_h_l1845_c7_9f69_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1845_c7_9f69]
signal n8_MUX_uxn_opcodes_h_l1845_c7_9f69_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1845_c7_9f69]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1845_c7_9f69]
signal result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1845_c7_9f69]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1845_c7_9f69]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1845_c7_9f69]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1848_c11_4775]
signal BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1848_c7_b999]
signal t8_MUX_uxn_opcodes_h_l1848_c7_b999_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1848_c7_b999_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1848_c7_b999]
signal n8_MUX_uxn_opcodes_h_l1848_c7_b999_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1848_c7_b999_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1848_c7_b999]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1848_c7_b999]
signal result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1848_c7_b999]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1848_c7_b999]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1848_c7_b999]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1851_c11_f831]
signal BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1851_c7_f68f]
signal n8_MUX_uxn_opcodes_h_l1851_c7_f68f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1851_c7_f68f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1851_c7_f68f]
signal result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1851_c7_f68f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1851_c7_f68f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1851_c7_f68f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1853_c30_9679]
signal sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_return_output : signed(3 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1856_c21_8e90]
signal BIN_OP_GT_uxn_opcodes_h_l1856_c21_8e90_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1856_c21_8e90_right : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1856_c21_8e90_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1856_c21_daa0]
signal MUX_uxn_opcodes_h_l1856_c21_daa0_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1856_c21_daa0_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1856_c21_daa0_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1856_c21_daa0_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_84a2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_vram_write := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_pc_updated := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb
BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_left,
BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_right,
BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_return_output);

-- t8_MUX_uxn_opcodes_h_l1832_c2_0399
t8_MUX_uxn_opcodes_h_l1832_c2_0399 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1832_c2_0399_cond,
t8_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue,
t8_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse,
t8_MUX_uxn_opcodes_h_l1832_c2_0399_return_output);

-- n8_MUX_uxn_opcodes_h_l1832_c2_0399
n8_MUX_uxn_opcodes_h_l1832_c2_0399 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1832_c2_0399_cond,
n8_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue,
n8_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse,
n8_MUX_uxn_opcodes_h_l1832_c2_0399_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399
result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399
result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399
result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399
result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399
result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399
result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_cond,
result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399
result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c
BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_left,
BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_right,
BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_return_output);

-- t8_MUX_uxn_opcodes_h_l1845_c7_9f69
t8_MUX_uxn_opcodes_h_l1845_c7_9f69 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1845_c7_9f69_cond,
t8_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue,
t8_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse,
t8_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output);

-- n8_MUX_uxn_opcodes_h_l1845_c7_9f69
n8_MUX_uxn_opcodes_h_l1845_c7_9f69 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1845_c7_9f69_cond,
n8_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue,
n8_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse,
n8_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69
result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69
result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_cond,
result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69
result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69
result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775
BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_left,
BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_right,
BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_return_output);

-- t8_MUX_uxn_opcodes_h_l1848_c7_b999
t8_MUX_uxn_opcodes_h_l1848_c7_b999 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1848_c7_b999_cond,
t8_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue,
t8_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse,
t8_MUX_uxn_opcodes_h_l1848_c7_b999_return_output);

-- n8_MUX_uxn_opcodes_h_l1848_c7_b999
n8_MUX_uxn_opcodes_h_l1848_c7_b999 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1848_c7_b999_cond,
n8_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue,
n8_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse,
n8_MUX_uxn_opcodes_h_l1848_c7_b999_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999
result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999
result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_cond,
result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999
result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999
result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831
BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831_left,
BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831_right,
BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831_return_output);

-- n8_MUX_uxn_opcodes_h_l1851_c7_f68f
n8_MUX_uxn_opcodes_h_l1851_c7_f68f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1851_c7_f68f_cond,
n8_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue,
n8_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse,
n8_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f
result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f
result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f
result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1853_c30_9679
sp_relative_shift_uxn_opcodes_h_l1853_c30_9679 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_ins,
sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_x,
sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_y,
sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1856_c21_8e90
BIN_OP_GT_uxn_opcodes_h_l1856_c21_8e90 : entity work.BIN_OP_GT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1856_c21_8e90_left,
BIN_OP_GT_uxn_opcodes_h_l1856_c21_8e90_right,
BIN_OP_GT_uxn_opcodes_h_l1856_c21_8e90_return_output);

-- MUX_uxn_opcodes_h_l1856_c21_daa0
MUX_uxn_opcodes_h_l1856_c21_daa0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1856_c21_daa0_cond,
MUX_uxn_opcodes_h_l1856_c21_daa0_iftrue,
MUX_uxn_opcodes_h_l1856_c21_daa0_iffalse,
MUX_uxn_opcodes_h_l1856_c21_daa0_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_return_output,
 t8_MUX_uxn_opcodes_h_l1832_c2_0399_return_output,
 n8_MUX_uxn_opcodes_h_l1832_c2_0399_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_return_output,
 t8_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output,
 n8_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_return_output,
 t8_MUX_uxn_opcodes_h_l1848_c7_b999_return_output,
 n8_MUX_uxn_opcodes_h_l1848_c7_b999_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831_return_output,
 n8_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output,
 sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1856_c21_8e90_return_output,
 MUX_uxn_opcodes_h_l1856_c21_daa0_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1832_c2_0399_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1832_c2_0399_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1832_c2_0399_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1832_c2_0399_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1832_c2_0399_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1832_c2_0399_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1837_c3_6c6b : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1832_c2_0399_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1842_c3_bb5c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1832_c2_0399_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1848_c7_b999_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1845_c7_9f69_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1848_c7_b999_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1845_c7_9f69_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1846_c3_6a7c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1848_c7_b999_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1848_c7_b999_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1851_c7_f68f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1855_c3_7604 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1856_c21_daa0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1856_c21_8e90_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1856_c21_8e90_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1856_c21_8e90_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1856_c21_daa0_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1856_c21_daa0_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1856_c21_daa0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1832_l1851_l1845_l1848_DUPLICATE_a65b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1851_l1845_l1848_DUPLICATE_ba07_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1851_l1845_l1848_DUPLICATE_0a85_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1851_l1845_l1848_DUPLICATE_167b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1851_l1848_DUPLICATE_624b_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1860_l1828_DUPLICATE_d8cb_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1837_c3_6c6b := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1837_c3_6c6b;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_MUX_uxn_opcodes_h_l1856_c21_daa0_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1846_c3_6a7c := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1846_c3_6a7c;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1855_c3_7604 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1855_c3_7604;
     VAR_MUX_uxn_opcodes_h_l1856_c21_daa0_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1842_c3_bb5c := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1842_c3_bb5c;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_right := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831_left := VAR_phase;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1856_c21_8e90_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1856_c21_8e90_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse := t8;
     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1832_c2_0399] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1832_c2_0399_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l1848_c11_4775] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_left;
     BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_return_output := BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1832_l1851_l1845_l1848_DUPLICATE_a65b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1832_l1851_l1845_l1848_DUPLICATE_a65b_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1832_c6_9abb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_left;
     BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_return_output := BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1832_c2_0399] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1832_c2_0399_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1851_l1845_l1848_DUPLICATE_167b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1851_l1845_l1848_DUPLICATE_167b_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1851_l1848_DUPLICATE_624b LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1851_l1848_DUPLICATE_624b_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1851_c11_f831] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831_left;
     BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831_return_output := BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l1856_c21_8e90] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1856_c21_8e90_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1856_c21_8e90_left;
     BIN_OP_GT_uxn_opcodes_h_l1856_c21_8e90_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1856_c21_8e90_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1856_c21_8e90_return_output := BIN_OP_GT_uxn_opcodes_h_l1856_c21_8e90_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1851_l1845_l1848_DUPLICATE_0a85 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1851_l1845_l1848_DUPLICATE_0a85_return_output := result.sp_relative_shift;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1832_c2_0399] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1832_c2_0399_return_output := result.is_pc_updated;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1832_c2_0399] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1832_c2_0399_return_output := result.is_vram_write;

     -- sp_relative_shift[uxn_opcodes_h_l1853_c30_9679] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_ins;
     sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_x;
     sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_return_output := sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1851_l1845_l1848_DUPLICATE_ba07 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1851_l1845_l1848_DUPLICATE_ba07_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1845_c11_726c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1832_c2_0399_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1832_c2_0399_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1832_c6_9abb_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1845_c7_9f69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1845_c7_9f69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_726c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1848_c7_b999_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1848_c7_b999_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1848_c11_4775_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1851_c7_f68f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1851_c11_f831_return_output;
     VAR_MUX_uxn_opcodes_h_l1856_c21_daa0_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1856_c21_8e90_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1851_l1845_l1848_DUPLICATE_0a85_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1851_l1845_l1848_DUPLICATE_0a85_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1851_l1845_l1848_DUPLICATE_0a85_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1851_l1845_l1848_DUPLICATE_ba07_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1851_l1845_l1848_DUPLICATE_ba07_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1851_l1845_l1848_DUPLICATE_ba07_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1851_l1845_l1848_DUPLICATE_167b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1851_l1845_l1848_DUPLICATE_167b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1851_l1845_l1848_DUPLICATE_167b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1851_l1848_DUPLICATE_624b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1851_l1848_DUPLICATE_624b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1832_l1851_l1845_l1848_DUPLICATE_a65b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1832_l1851_l1845_l1848_DUPLICATE_a65b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1832_l1851_l1845_l1848_DUPLICATE_a65b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1832_l1851_l1845_l1848_DUPLICATE_a65b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1832_c2_0399_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1832_c2_0399_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1832_c2_0399_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1832_c2_0399_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1853_c30_9679_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1832_c2_0399] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1832_c2_0399] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1851_c7_f68f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1851_c7_f68f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1851_c7_f68f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1832_c2_0399] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1851_c7_f68f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output;

     -- n8_MUX[uxn_opcodes_h_l1851_c7_f68f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1851_c7_f68f_cond <= VAR_n8_MUX_uxn_opcodes_h_l1851_c7_f68f_cond;
     n8_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue;
     n8_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output := n8_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output;

     -- MUX[uxn_opcodes_h_l1856_c21_daa0] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1856_c21_daa0_cond <= VAR_MUX_uxn_opcodes_h_l1856_c21_daa0_cond;
     MUX_uxn_opcodes_h_l1856_c21_daa0_iftrue <= VAR_MUX_uxn_opcodes_h_l1856_c21_daa0_iftrue;
     MUX_uxn_opcodes_h_l1856_c21_daa0_iffalse <= VAR_MUX_uxn_opcodes_h_l1856_c21_daa0_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1856_c21_daa0_return_output := MUX_uxn_opcodes_h_l1856_c21_daa0_return_output;

     -- t8_MUX[uxn_opcodes_h_l1848_c7_b999] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1848_c7_b999_cond <= VAR_t8_MUX_uxn_opcodes_h_l1848_c7_b999_cond;
     t8_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue;
     t8_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1848_c7_b999_return_output := t8_MUX_uxn_opcodes_h_l1848_c7_b999_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1832_c2_0399] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue := VAR_MUX_uxn_opcodes_h_l1856_c21_daa0_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1848_c7_b999_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1848_c7_b999] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1848_c7_b999] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1848_c7_b999] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_return_output;

     -- n8_MUX[uxn_opcodes_h_l1848_c7_b999] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1848_c7_b999_cond <= VAR_n8_MUX_uxn_opcodes_h_l1848_c7_b999_cond;
     n8_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue;
     n8_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1848_c7_b999_return_output := n8_MUX_uxn_opcodes_h_l1848_c7_b999_return_output;

     -- t8_MUX[uxn_opcodes_h_l1845_c7_9f69] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1845_c7_9f69_cond <= VAR_t8_MUX_uxn_opcodes_h_l1845_c7_9f69_cond;
     t8_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue;
     t8_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output := t8_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1851_c7_f68f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1848_c7_b999] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1848_c7_b999_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1848_c7_b999_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1848_c7_b999_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1848_c7_b999_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1848_c7_b999_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1851_c7_f68f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1845_c7_9f69] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output;

     -- t8_MUX[uxn_opcodes_h_l1832_c2_0399] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1832_c2_0399_cond <= VAR_t8_MUX_uxn_opcodes_h_l1832_c2_0399_cond;
     t8_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue;
     t8_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1832_c2_0399_return_output := t8_MUX_uxn_opcodes_h_l1832_c2_0399_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1845_c7_9f69] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1845_c7_9f69] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1845_c7_9f69] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1848_c7_b999] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_return_output := result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_return_output;

     -- n8_MUX[uxn_opcodes_h_l1845_c7_9f69] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1845_c7_9f69_cond <= VAR_n8_MUX_uxn_opcodes_h_l1845_c7_9f69_cond;
     n8_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue;
     n8_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output := n8_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1848_c7_b999_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1832_c2_0399_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1832_c2_0399] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1832_c2_0399] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1845_c7_9f69] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output := result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1832_c2_0399] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_return_output;

     -- n8_MUX[uxn_opcodes_h_l1832_c2_0399] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1832_c2_0399_cond <= VAR_n8_MUX_uxn_opcodes_h_l1832_c2_0399_cond;
     n8_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue;
     n8_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1832_c2_0399_return_output := n8_MUX_uxn_opcodes_h_l1832_c2_0399_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1832_c2_0399] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1832_c2_0399_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_9f69_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1832_c2_0399] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_return_output := result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1860_l1828_DUPLICATE_d8cb LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1860_l1828_DUPLICATE_d8cb_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_84a2(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1832_c2_0399_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1832_c2_0399_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1832_c2_0399_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1832_c2_0399_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1832_c2_0399_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1832_c2_0399_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1832_c2_0399_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1832_c2_0399_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1832_c2_0399_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1860_l1828_DUPLICATE_d8cb_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1860_l1828_DUPLICATE_d8cb_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
