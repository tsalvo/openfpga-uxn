-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 48
entity dei_0CLK_fcb212cd is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_device_ram_read : in unsigned(15 downto 0);
 return_output : out opcode_result_t);
end dei_0CLK_fcb212cd;
architecture arch of dei_0CLK_fcb212cd is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal has_written_to_t : unsigned(0 downto 0) := to_unsigned(0, 1);
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal device_in_result : device_in_result_t := device_in_result_t_NULL;
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_has_written_to_t : unsigned(0 downto 0);
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_device_in_result : device_in_result_t;
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l380_c6_6417]
signal BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l391_c7_9e2d]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output : unsigned(0 downto 0);

-- device_in_result_MUX[uxn_opcodes_h_l380_c2_1e0d]
signal device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_cond : unsigned(0 downto 0);
signal device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output : device_in_result_t;

-- result_is_device_ram_16bit_MUX[uxn_opcodes_h_l380_c2_1e0d]
signal result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_cond : unsigned(0 downto 0);
signal result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output : unsigned(0 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l380_c2_1e0d]
signal result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l380_c2_1e0d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output : unsigned(0 downto 0);

-- result_is_device_ram_write_MUX[uxn_opcodes_h_l380_c2_1e0d]
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_cond : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l380_c2_1e0d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l380_c2_1e0d]
signal result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l380_c2_1e0d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l380_c2_1e0d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l380_c2_1e0d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l380_c2_1e0d]
signal t8_MUX_uxn_opcodes_h_l380_c2_1e0d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output : unsigned(7 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l380_c2_1e0d]
signal has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l391_c11_595b]
signal BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l395_c1_b803]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_return_output : unsigned(0 downto 0);

-- device_in_result_MUX[uxn_opcodes_h_l391_c7_9e2d]
signal device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_cond : unsigned(0 downto 0);
signal device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output : device_in_result_t;

-- result_device_ram_address_MUX[uxn_opcodes_h_l391_c7_9e2d]
signal result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l391_c7_9e2d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l391_c7_9e2d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l391_c7_9e2d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l391_c7_9e2d]
signal result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l391_c7_9e2d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l391_c7_9e2d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l391_c7_9e2d]
signal t8_MUX_uxn_opcodes_h_l391_c7_9e2d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output : unsigned(7 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l391_c7_9e2d]
signal has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l393_c30_0d84]
signal sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l397_c9_c763]
signal BIN_OP_EQ_uxn_opcodes_h_l397_c9_c763_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l397_c9_c763_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l397_c9_c763_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l397_c9_3c9d]
signal MUX_uxn_opcodes_h_l397_c9_3c9d_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l397_c9_3c9d_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l397_c9_3c9d_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l397_c9_3c9d_return_output : unsigned(7 downto 0);

-- UNARY_OP_NOT[uxn_opcodes_h_l398_c8_e9ea]
signal UNARY_OP_NOT_uxn_opcodes_h_l398_c8_e9ea_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_uxn_opcodes_h_l398_c8_e9ea_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l398_c1_75e1]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_return_output : unsigned(0 downto 0);

-- device_in_result_MUX[uxn_opcodes_h_l398_c3_481c]
signal device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_cond : unsigned(0 downto 0);
signal device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_iftrue : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_iffalse : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_return_output : device_in_result_t;

-- result_device_ram_address_MUX[uxn_opcodes_h_l398_c3_481c]
signal result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l398_c3_481c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l398_c3_481c]
signal result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l398_c3_481c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l398_c3_481c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_return_output : unsigned(3 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l398_c3_481c]
signal has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_return_output : unsigned(0 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_h_l399_c37_33fc]
signal BIN_OP_MINUS_uxn_opcodes_h_l399_c37_33fc_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l399_c37_33fc_right : unsigned(1 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l399_c37_33fc_return_output : unsigned(7 downto 0);

-- device_in[uxn_opcodes_h_l399_c23_8777]
signal device_in_uxn_opcodes_h_l399_c23_8777_CLOCK_ENABLE : unsigned(0 downto 0);
signal device_in_uxn_opcodes_h_l399_c23_8777_device_address : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l399_c23_8777_phase : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l399_c23_8777_previous_device_ram_read : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l399_c23_8777_return_output : device_in_result_t;

-- UNARY_OP_NOT[uxn_opcodes_h_l402_c9_e47d]
signal UNARY_OP_NOT_uxn_opcodes_h_l402_c9_e47d_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_uxn_opcodes_h_l402_c9_e47d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l402_c4_214f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l402_c4_214f]
signal result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l402_c4_214f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l402_c4_214f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_return_output : unsigned(3 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l402_c4_214f]
signal has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_return_output : unsigned(0 downto 0);

function CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6( ref_toks_0 : device_in_result_t;
 ref_toks_1 : unsigned) return device_in_result_t is
 
  variable base : device_in_result_t; 
  variable return_output : device_in_result_t;
begin
      base := ref_toks_0;
      base.is_dei_done := ref_toks_1;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_8a80( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_device_ram_16bit := ref_toks_1;
      base.device_ram_address := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_device_ram_write := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.u8_value := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_sp_shift := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417
BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_left,
BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_right,
BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output);

-- device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d
device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_cond,
device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue,
device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse,
device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output);

-- result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d
result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_cond,
result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue,
result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse,
result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d
result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d
result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output);

-- result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d
result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_cond,
result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue,
result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse,
result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d
result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d
result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_cond,
result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d
result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d
result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output);

-- t8_MUX_uxn_opcodes_h_l380_c2_1e0d
t8_MUX_uxn_opcodes_h_l380_c2_1e0d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l380_c2_1e0d_cond,
t8_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue,
t8_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse,
t8_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d
has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_cond,
has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b
BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_left,
BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_right,
BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_return_output);

-- device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d
device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_cond,
device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue,
device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse,
device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d
result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d
result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d
result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d
result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_cond,
result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d
result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d
result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output);

-- t8_MUX_uxn_opcodes_h_l391_c7_9e2d
t8_MUX_uxn_opcodes_h_l391_c7_9e2d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l391_c7_9e2d_cond,
t8_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue,
t8_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse,
t8_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d
has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_cond,
has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output);

-- sp_relative_shift_uxn_opcodes_h_l393_c30_0d84
sp_relative_shift_uxn_opcodes_h_l393_c30_0d84 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_ins,
sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_x,
sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_y,
sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l397_c9_c763
BIN_OP_EQ_uxn_opcodes_h_l397_c9_c763 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l397_c9_c763_left,
BIN_OP_EQ_uxn_opcodes_h_l397_c9_c763_right,
BIN_OP_EQ_uxn_opcodes_h_l397_c9_c763_return_output);

-- MUX_uxn_opcodes_h_l397_c9_3c9d
MUX_uxn_opcodes_h_l397_c9_3c9d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l397_c9_3c9d_cond,
MUX_uxn_opcodes_h_l397_c9_3c9d_iftrue,
MUX_uxn_opcodes_h_l397_c9_3c9d_iffalse,
MUX_uxn_opcodes_h_l397_c9_3c9d_return_output);

-- UNARY_OP_NOT_uxn_opcodes_h_l398_c8_e9ea
UNARY_OP_NOT_uxn_opcodes_h_l398_c8_e9ea : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_uxn_opcodes_h_l398_c8_e9ea_expr,
UNARY_OP_NOT_uxn_opcodes_h_l398_c8_e9ea_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_return_output);

-- device_in_result_MUX_uxn_opcodes_h_l398_c3_481c
device_in_result_MUX_uxn_opcodes_h_l398_c3_481c : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_cond,
device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_iftrue,
device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_iffalse,
device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c
result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c
result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c
result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_cond,
result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c
result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c
has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_cond,
has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l399_c37_33fc
BIN_OP_MINUS_uxn_opcodes_h_l399_c37_33fc : entity work.BIN_OP_MINUS_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l399_c37_33fc_left,
BIN_OP_MINUS_uxn_opcodes_h_l399_c37_33fc_right,
BIN_OP_MINUS_uxn_opcodes_h_l399_c37_33fc_return_output);

-- device_in_uxn_opcodes_h_l399_c23_8777
device_in_uxn_opcodes_h_l399_c23_8777 : entity work.device_in_0CLK_85463cfa port map (
clk,
device_in_uxn_opcodes_h_l399_c23_8777_CLOCK_ENABLE,
device_in_uxn_opcodes_h_l399_c23_8777_device_address,
device_in_uxn_opcodes_h_l399_c23_8777_phase,
device_in_uxn_opcodes_h_l399_c23_8777_previous_device_ram_read,
device_in_uxn_opcodes_h_l399_c23_8777_return_output);

-- UNARY_OP_NOT_uxn_opcodes_h_l402_c9_e47d
UNARY_OP_NOT_uxn_opcodes_h_l402_c9_e47d : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_uxn_opcodes_h_l402_c9_e47d_expr,
UNARY_OP_NOT_uxn_opcodes_h_l402_c9_e47d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f
result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f
result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_cond,
result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f
result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f
has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_cond,
has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_device_ram_read,
 -- Registers
 has_written_to_t,
 t8,
 device_in_result,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output,
 device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output,
 result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output,
 result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output,
 t8_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_return_output,
 device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output,
 t8_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output,
 sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l397_c9_c763_return_output,
 MUX_uxn_opcodes_h_l397_c9_3c9d_return_output,
 UNARY_OP_NOT_uxn_opcodes_h_l398_c8_e9ea_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_return_output,
 device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l399_c37_33fc_return_output,
 device_in_uxn_opcodes_h_l399_c23_8777_return_output,
 UNARY_OP_NOT_uxn_opcodes_h_l402_c9_e47d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_device_ram_read : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse : unsigned(0 downto 0);
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue : device_in_result_t;
 variable VAR_device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6_uxn_opcodes_h_l380_c2_1e0d_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_cond : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_16bit_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_16bit_d41d_uxn_opcodes_h_l380_c2_1e0d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_cond : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l380_c2_1e0d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l385_c3_4ba5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_TRUE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l380_c2_1e0d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l380_c2_1e0d_cond : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_iffalse : unsigned(0 downto 0);
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l391_c7_9e2d_cond : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l397_c9_3c9d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l397_c9_c763_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l397_c9_c763_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l397_c9_c763_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l397_c9_3c9d_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l397_c9_3c9d_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l397_c9_3c9d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d_uxn_opcodes_h_l398_c8_f79d_return_output : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l398_c8_e9ea_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l398_c8_e9ea_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_iffalse : unsigned(0 downto 0);
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_iftrue : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_iffalse : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_cond : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_cond : unsigned(0 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l399_c23_8777_device_address : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l399_c23_8777_phase : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l399_c23_8777_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l399_c37_33fc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l399_c37_33fc_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l399_c37_33fc_return_output : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l399_c23_8777_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l399_c23_8777_return_output : device_in_result_t;
 variable VAR_CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d_uxn_opcodes_h_l400_c32_3b36_return_output : unsigned(7 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l402_c9_e47d_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l402_c9_e47d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l404_c5_01f6 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_cond : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d_uxn_opcodes_h_l405_c23_2986_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l380_l391_l398_DUPLICATE_19c6_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l380_l391_l398_DUPLICATE_3112_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l380_l402_l391_l398_DUPLICATE_1d93_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l380_l391_DUPLICATE_d8d7_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l402_l391_l398_DUPLICATE_6465_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l402_l391_l398_DUPLICATE_7e17_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8a80_uxn_opcodes_h_l414_l374_DUPLICATE_9223_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_has_written_to_t : unsigned(0 downto 0);
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_device_in_result : device_in_result_t;
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_has_written_to_t := has_written_to_t;
  REG_VAR_t8 := t8;
  REG_VAR_device_in_result := device_in_result;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_right := to_unsigned(0, 1);
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_iffalse := to_unsigned(0, 1);
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l399_c37_33fc_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l404_c5_01f6 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l404_c5_01f6;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_iffalse := to_unsigned(1, 1);
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_iftrue := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_right := to_unsigned(1, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_iftrue := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l397_c9_c763_right := to_unsigned(2, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l385_c3_4ba5 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l385_c3_4ba5;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_device_ram_read := previous_device_ram_read;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse := VAR_CLOCK_ENABLE;
     VAR_device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue := device_in_result;
     VAR_device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_iffalse := device_in_result;
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l402_c9_e47d_expr := has_written_to_t;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue := has_written_to_t;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_iftrue := has_written_to_t;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_iffalse := has_written_to_t;
     VAR_sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l397_c9_c763_left := VAR_phase;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l399_c37_33fc_left := VAR_phase;
     VAR_device_in_uxn_opcodes_h_l399_c23_8777_previous_device_ram_read := resize(VAR_previous_device_ram_read, 8);
     VAR_MUX_uxn_opcodes_h_l397_c9_3c9d_iftrue := VAR_previous_stack_read;
     VAR_MUX_uxn_opcodes_h_l397_c9_3c9d_iffalse := t8;
     VAR_t8_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue := t8;
     -- UNARY_OP_NOT[uxn_opcodes_h_l402_c9_e47d] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_uxn_opcodes_h_l402_c9_e47d_expr <= VAR_UNARY_OP_NOT_uxn_opcodes_h_l402_c9_e47d_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l402_c9_e47d_return_output := UNARY_OP_NOT_uxn_opcodes_h_l402_c9_e47d_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l402_l391_l398_DUPLICATE_7e17 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l402_l391_l398_DUPLICATE_7e17_return_output := result.is_opc_done;

     -- result_is_device_ram_16bit_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_16bit_d41d[uxn_opcodes_h_l380_c2_1e0d] LATENCY=0
     VAR_result_is_device_ram_16bit_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_16bit_d41d_uxn_opcodes_h_l380_c2_1e0d_return_output := result.is_device_ram_16bit;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l402_l391_l398_DUPLICATE_6465 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l402_l391_l398_DUPLICATE_6465_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d[uxn_opcodes_h_l405_c23_2986] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d_uxn_opcodes_h_l405_c23_2986_return_output := device_in_result.dei_value;

     -- CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l380_l391_l398_DUPLICATE_19c6 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l380_l391_l398_DUPLICATE_19c6_return_output := result.device_ram_address;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l380_l402_l391_l398_DUPLICATE_1d93 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l380_l402_l391_l398_DUPLICATE_1d93_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l391_c11_595b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_left;
     BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_return_output := BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_return_output;

     -- result_is_sp_shift_TRUE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d[uxn_opcodes_h_l380_c2_1e0d] LATENCY=0
     VAR_result_is_sp_shift_TRUE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l380_c2_1e0d_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l397_c9_c763] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l397_c9_c763_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l397_c9_c763_left;
     BIN_OP_EQ_uxn_opcodes_h_l397_c9_c763_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l397_c9_c763_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l397_c9_c763_return_output := BIN_OP_EQ_uxn_opcodes_h_l397_c9_c763_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l380_l391_DUPLICATE_d8d7 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l380_l391_DUPLICATE_d8d7_return_output := result.sp_relative_shift;

     -- BIN_OP_MINUS[uxn_opcodes_h_l399_c37_33fc] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l399_c37_33fc_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l399_c37_33fc_left;
     BIN_OP_MINUS_uxn_opcodes_h_l399_c37_33fc_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l399_c37_33fc_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l399_c37_33fc_return_output := BIN_OP_MINUS_uxn_opcodes_h_l399_c37_33fc_return_output;

     -- result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d[uxn_opcodes_h_l380_c2_1e0d] LATENCY=0
     VAR_result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l380_c2_1e0d_return_output := result.is_device_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l380_l391_l398_DUPLICATE_3112 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l380_l391_l398_DUPLICATE_3112_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l380_c6_6417] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_left;
     BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_return_output := BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_return_output;

     -- CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d[uxn_opcodes_h_l398_c8_f79d] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d_uxn_opcodes_h_l398_c8_f79d_return_output := device_in_result.is_dei_done;

     -- sp_relative_shift[uxn_opcodes_h_l393_c30_0d84] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_ins;
     sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_x <= VAR_sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_x;
     sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_y <= VAR_sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_return_output := sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_return_output;

     -- device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6[uxn_opcodes_h_l380_c2_1e0d] LATENCY=0
     VAR_device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6_uxn_opcodes_h_l380_c2_1e0d_return_output := CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6(
     device_in_result,
     to_unsigned(0, 1));

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_return_output;
     VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l380_c2_1e0d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l380_c6_6417_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l391_c7_9e2d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l391_c11_595b_return_output;
     VAR_MUX_uxn_opcodes_h_l397_c9_3c9d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l397_c9_c763_return_output;
     VAR_device_in_uxn_opcodes_h_l399_c23_8777_phase := VAR_BIN_OP_MINUS_uxn_opcodes_h_l399_c37_33fc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l380_l391_DUPLICATE_d8d7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l380_l391_DUPLICATE_d8d7_return_output;
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l398_c8_e9ea_expr := VAR_CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d_uxn_opcodes_h_l398_c8_f79d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l402_l391_l398_DUPLICATE_7e17_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l402_l391_l398_DUPLICATE_7e17_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l402_l391_l398_DUPLICATE_7e17_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l380_l391_l398_DUPLICATE_3112_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l380_l391_l398_DUPLICATE_3112_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l380_l391_l398_DUPLICATE_3112_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l402_l391_l398_DUPLICATE_6465_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l402_l391_l398_DUPLICATE_6465_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l402_l391_l398_DUPLICATE_6465_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_iftrue := VAR_CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d_uxn_opcodes_h_l405_c23_2986_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l380_l391_l398_DUPLICATE_19c6_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l380_l391_l398_DUPLICATE_19c6_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l380_l391_l398_DUPLICATE_19c6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l380_l402_l391_l398_DUPLICATE_1d93_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l380_l402_l391_l398_DUPLICATE_1d93_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l380_l402_l391_l398_DUPLICATE_1d93_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l380_l402_l391_l398_DUPLICATE_1d93_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l402_c9_e47d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l402_c9_e47d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l402_c9_e47d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l402_c9_e47d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l402_c9_e47d_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue := VAR_device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6_uxn_opcodes_h_l380_c2_1e0d_return_output;
     VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse := VAR_result_is_device_ram_16bit_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_16bit_d41d_uxn_opcodes_h_l380_c2_1e0d_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse := VAR_result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l380_c2_1e0d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue := VAR_result_is_sp_shift_TRUE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l380_c2_1e0d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l393_c30_0d84_return_output;
     -- MUX[uxn_opcodes_h_l397_c9_3c9d] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l397_c9_3c9d_cond <= VAR_MUX_uxn_opcodes_h_l397_c9_3c9d_cond;
     MUX_uxn_opcodes_h_l397_c9_3c9d_iftrue <= VAR_MUX_uxn_opcodes_h_l397_c9_3c9d_iftrue;
     MUX_uxn_opcodes_h_l397_c9_3c9d_iffalse <= VAR_MUX_uxn_opcodes_h_l397_c9_3c9d_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l397_c9_3c9d_return_output := MUX_uxn_opcodes_h_l397_c9_3c9d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l402_c4_214f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_return_output;

     -- result_is_device_ram_write_MUX[uxn_opcodes_h_l380_c2_1e0d] LATENCY=0
     -- Inputs
     result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_cond <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_cond;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse;
     -- Outputs
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output := result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output;

     -- UNARY_OP_NOT[uxn_opcodes_h_l398_c8_e9ea] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_uxn_opcodes_h_l398_c8_e9ea_expr <= VAR_UNARY_OP_NOT_uxn_opcodes_h_l398_c8_e9ea_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l398_c8_e9ea_return_output := UNARY_OP_NOT_uxn_opcodes_h_l398_c8_e9ea_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l391_c7_9e2d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output;

     -- result_is_device_ram_16bit_MUX[uxn_opcodes_h_l380_c2_1e0d] LATENCY=0
     -- Inputs
     result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_cond <= VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_cond;
     result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue <= VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue;
     result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse <= VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse;
     -- Outputs
     VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output := result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l402_c4_214f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l402_c4_214f] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_return_output := has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l402_c4_214f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l402_c4_214f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_return_output := result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l391_c7_9e2d] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l391_c7_9e2d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output;
     VAR_device_in_uxn_opcodes_h_l399_c23_8777_device_address := VAR_MUX_uxn_opcodes_h_l397_c9_3c9d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse := VAR_MUX_uxn_opcodes_h_l397_c9_3c9d_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l398_c8_e9ea_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l398_c8_e9ea_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l398_c8_e9ea_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l398_c8_e9ea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l398_c8_e9ea_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l398_c8_e9ea_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l398_c8_e9ea_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l398_c8_e9ea_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_iffalse := VAR_has_written_to_t_MUX_uxn_opcodes_h_l402_c4_214f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l402_c4_214f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l402_c4_214f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l402_c4_214f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l402_c4_214f_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l380_c2_1e0d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l398_c3_481c] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_return_output := has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l398_c3_481c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l380_c2_1e0d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l398_c3_481c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_return_output := result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l395_c1_b803] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l398_c3_481c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_return_output;

     -- t8_MUX[uxn_opcodes_h_l391_c7_9e2d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l391_c7_9e2d_cond <= VAR_t8_MUX_uxn_opcodes_h_l391_c7_9e2d_cond;
     t8_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue;
     t8_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output := t8_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l398_c3_481c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_return_output;

     -- Submodule level 3
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l395_c1_b803_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse := VAR_has_written_to_t_MUX_uxn_opcodes_h_l398_c3_481c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l398_c3_481c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l398_c3_481c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l398_c3_481c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l398_c3_481c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse := VAR_t8_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l391_c7_9e2d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output := result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l391_c7_9e2d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l391_c7_9e2d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l391_c7_9e2d] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output := has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l398_c1_75e1] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l391_c7_9e2d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output;

     -- t8_MUX[uxn_opcodes_h_l380_c2_1e0d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l380_c2_1e0d_cond <= VAR_t8_MUX_uxn_opcodes_h_l380_c2_1e0d_cond;
     t8_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue;
     t8_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output := t8_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output;

     -- Submodule level 4
     VAR_device_in_uxn_opcodes_h_l399_c23_8777_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l398_c1_75e1_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse := VAR_has_written_to_t_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l380_c2_1e0d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l380_c2_1e0d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l380_c2_1e0d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output := result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l380_c2_1e0d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output;

     -- device_in[uxn_opcodes_h_l399_c23_8777] LATENCY=0
     -- Clock enable
     device_in_uxn_opcodes_h_l399_c23_8777_CLOCK_ENABLE <= VAR_device_in_uxn_opcodes_h_l399_c23_8777_CLOCK_ENABLE;
     -- Inputs
     device_in_uxn_opcodes_h_l399_c23_8777_device_address <= VAR_device_in_uxn_opcodes_h_l399_c23_8777_device_address;
     device_in_uxn_opcodes_h_l399_c23_8777_phase <= VAR_device_in_uxn_opcodes_h_l399_c23_8777_phase;
     device_in_uxn_opcodes_h_l399_c23_8777_previous_device_ram_read <= VAR_device_in_uxn_opcodes_h_l399_c23_8777_previous_device_ram_read;
     -- Outputs
     VAR_device_in_uxn_opcodes_h_l399_c23_8777_return_output := device_in_uxn_opcodes_h_l399_c23_8777_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l380_c2_1e0d] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output := has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output;

     -- Submodule level 5
     VAR_device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_iftrue := VAR_device_in_uxn_opcodes_h_l399_c23_8777_return_output;
     REG_VAR_has_written_to_t := VAR_has_written_to_t_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output;
     -- CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d[uxn_opcodes_h_l400_c32_3b36] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d_uxn_opcodes_h_l400_c32_3b36_return_output := VAR_device_in_uxn_opcodes_h_l399_c23_8777_return_output.device_ram_address;

     -- device_in_result_MUX[uxn_opcodes_h_l398_c3_481c] LATENCY=0
     -- Inputs
     device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_cond <= VAR_device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_cond;
     device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_iftrue <= VAR_device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_iftrue;
     device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_iffalse <= VAR_device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_iffalse;
     -- Outputs
     VAR_device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_return_output := device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_return_output;

     -- Submodule level 6
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_iftrue := VAR_CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d_uxn_opcodes_h_l400_c32_3b36_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse := VAR_device_in_result_MUX_uxn_opcodes_h_l398_c3_481c_return_output;
     -- device_in_result_MUX[uxn_opcodes_h_l391_c7_9e2d] LATENCY=0
     -- Inputs
     device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_cond <= VAR_device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_cond;
     device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue <= VAR_device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue;
     device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse <= VAR_device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse;
     -- Outputs
     VAR_device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output := device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output;

     -- result_device_ram_address_MUX[uxn_opcodes_h_l398_c3_481c] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_return_output;

     -- Submodule level 7
     VAR_device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse := VAR_device_in_result_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l398_c3_481c_return_output;
     -- device_in_result_MUX[uxn_opcodes_h_l380_c2_1e0d] LATENCY=0
     -- Inputs
     device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_cond <= VAR_device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_cond;
     device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue <= VAR_device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue;
     device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse <= VAR_device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse;
     -- Outputs
     VAR_device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output := device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output;

     -- result_device_ram_address_MUX[uxn_opcodes_h_l391_c7_9e2d] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output;

     -- Submodule level 8
     REG_VAR_device_in_result := VAR_device_in_result_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l391_c7_9e2d_return_output;
     -- result_device_ram_address_MUX[uxn_opcodes_h_l380_c2_1e0d] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output;

     -- Submodule level 9
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8a80_uxn_opcodes_h_l414_l374_DUPLICATE_9223 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8a80_uxn_opcodes_h_l414_l374_DUPLICATE_9223_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8a80(
     result,
     VAR_result_is_device_ram_16bit_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output,
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output,
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l380_c2_1e0d_return_output);

     -- Submodule level 10
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8a80_uxn_opcodes_h_l414_l374_DUPLICATE_9223_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8a80_uxn_opcodes_h_l414_l374_DUPLICATE_9223_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_has_written_to_t <= REG_VAR_has_written_to_t;
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_device_in_result <= REG_VAR_device_in_result;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     has_written_to_t <= REG_COMB_has_written_to_t;
     t8 <= REG_COMB_t8;
     device_in_result <= REG_COMB_device_in_result;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
