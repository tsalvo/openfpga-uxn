-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 32
entity nip2_0CLK_b7103d16 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(15 downto 0);
 return_output : out opcode_result_t);
end nip2_0CLK_b7103d16;
architecture arch of nip2_0CLK_b7103d16 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1964_c6_ff97]
signal BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1964_c2_c167]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1964_c2_c167]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1964_c2_c167]
signal result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1964_c2_c167]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1964_c2_c167]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1964_c2_c167]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1964_c2_c167]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l1964_c2_c167]
signal t16_MUX_uxn_opcodes_h_l1964_c2_c167_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1964_c2_c167_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1972_c11_6cc2]
signal BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1972_c7_5c34]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1972_c7_5c34]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1972_c7_5c34]
signal result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1972_c7_5c34]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1972_c7_5c34]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1972_c7_5c34]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1972_c7_5c34]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l1972_c7_5c34]
signal t16_MUX_uxn_opcodes_h_l1972_c7_5c34_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1974_c30_998c]
signal sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1976_c11_e5d2]
signal BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1976_c7_b851]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1976_c7_b851]
signal result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1976_c7_b851]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1976_c7_b851]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1976_c7_b851]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1976_c7_b851]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_return_output : unsigned(3 downto 0);

-- t16_MUX[uxn_opcodes_h_l1976_c7_b851]
signal t16_MUX_uxn_opcodes_h_l1976_c7_b851_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1976_c7_b851_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1983_c11_6e6e]
signal BIN_OP_EQ_uxn_opcodes_h_l1983_c11_6e6e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1983_c11_6e6e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1983_c11_6e6e_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1983_c7_a875]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1983_c7_a875]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1983_c7_a875]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8152( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_stack_operation_16bit := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_stack_write := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97
BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_left,
BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_right,
BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167
result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167
result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_cond,
result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167
result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167
result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167
result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_return_output);

-- t16_MUX_uxn_opcodes_h_l1964_c2_c167
t16_MUX_uxn_opcodes_h_l1964_c2_c167 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1964_c2_c167_cond,
t16_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue,
t16_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse,
t16_MUX_uxn_opcodes_h_l1964_c2_c167_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2
BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_left,
BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_right,
BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34
result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34
result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_cond,
result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34
result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34
result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34
result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output);

-- t16_MUX_uxn_opcodes_h_l1972_c7_5c34
t16_MUX_uxn_opcodes_h_l1972_c7_5c34 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1972_c7_5c34_cond,
t16_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue,
t16_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse,
t16_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1974_c30_998c
sp_relative_shift_uxn_opcodes_h_l1974_c30_998c : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_ins,
sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_x,
sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_y,
sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2
BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_left,
BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_right,
BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851
result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851
result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_cond,
result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851
result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851
result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_return_output);

-- t16_MUX_uxn_opcodes_h_l1976_c7_b851
t16_MUX_uxn_opcodes_h_l1976_c7_b851 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1976_c7_b851_cond,
t16_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue,
t16_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse,
t16_MUX_uxn_opcodes_h_l1976_c7_b851_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1983_c11_6e6e
BIN_OP_EQ_uxn_opcodes_h_l1983_c11_6e6e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1983_c11_6e6e_left,
BIN_OP_EQ_uxn_opcodes_h_l1983_c11_6e6e_right,
BIN_OP_EQ_uxn_opcodes_h_l1983_c11_6e6e_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875
result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875
result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_return_output,
 t16_MUX_uxn_opcodes_h_l1964_c2_c167_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output,
 t16_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output,
 sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_return_output,
 t16_MUX_uxn_opcodes_h_l1976_c7_b851_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1983_c11_6e6e_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1969_c3_71c0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1964_c2_c167_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1964_c2_c167_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1976_c7_b851_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1972_c7_5c34_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1980_c3_adfc : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1976_c7_b851_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_6e6e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_6e6e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_6e6e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1976_l1964_DUPLICATE_7310_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1976_l1964_l1972_DUPLICATE_40fd_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1964_l1972_DUPLICATE_c5c9_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1964_l1983_l1972_DUPLICATE_0e48_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1976_l1972_DUPLICATE_e4f1_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1976_l1983_l1972_DUPLICATE_cbf0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1976_l1983_l1972_DUPLICATE_6898_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1989_l1960_DUPLICATE_9348_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1980_c3_adfc := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1980_c3_adfc;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1969_c3_71c0 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1969_c3_71c0;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_6e6e_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_y := resize(to_signed(-2, 3), 4);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_6e6e_left := VAR_phase;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue := VAR_previous_stack_read;
     VAR_t16_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue := VAR_previous_stack_read;
     VAR_t16_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse := t16;
     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1976_l1964_l1972_DUPLICATE_40fd LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1976_l1964_l1972_DUPLICATE_40fd_return_output := result.u16_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1976_l1964_DUPLICATE_7310 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1976_l1964_DUPLICATE_7310_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1976_c11_e5d2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_left;
     BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_return_output := BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1964_c6_ff97] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_left;
     BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_return_output := BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1974_c30_998c] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_ins;
     sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_x;
     sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_return_output := sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1964_l1972_DUPLICATE_c5c9 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1964_l1972_DUPLICATE_c5c9_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1976_l1983_l1972_DUPLICATE_6898 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1976_l1983_l1972_DUPLICATE_6898_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1983_c11_6e6e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1983_c11_6e6e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_6e6e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1983_c11_6e6e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_6e6e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_6e6e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1983_c11_6e6e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1972_c11_6cc2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_left;
     BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_return_output := BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1976_l1983_l1972_DUPLICATE_cbf0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1976_l1983_l1972_DUPLICATE_cbf0_return_output := result.is_stack_operation_16bit;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1976_l1972_DUPLICATE_e4f1 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1976_l1972_DUPLICATE_e4f1_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1964_l1983_l1972_DUPLICATE_0e48 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1964_l1983_l1972_DUPLICATE_0e48_return_output := result.is_stack_write;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1964_c2_c167_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c6_ff97_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1972_c7_5c34_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_6cc2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1976_c7_b851_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1976_c11_e5d2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_6e6e_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_6e6e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_6e6e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1964_l1972_DUPLICATE_c5c9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1964_l1972_DUPLICATE_c5c9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1976_l1964_l1972_DUPLICATE_40fd_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1976_l1964_l1972_DUPLICATE_40fd_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1976_l1964_l1972_DUPLICATE_40fd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1976_l1983_l1972_DUPLICATE_6898_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1976_l1983_l1972_DUPLICATE_6898_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1976_l1983_l1972_DUPLICATE_6898_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1976_l1964_DUPLICATE_7310_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1976_l1964_DUPLICATE_7310_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1976_l1983_l1972_DUPLICATE_cbf0_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1976_l1983_l1972_DUPLICATE_cbf0_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1976_l1983_l1972_DUPLICATE_cbf0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1964_l1983_l1972_DUPLICATE_0e48_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1964_l1983_l1972_DUPLICATE_0e48_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1964_l1983_l1972_DUPLICATE_0e48_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1976_l1972_DUPLICATE_e4f1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1976_l1972_DUPLICATE_e4f1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1974_c30_998c_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1983_c7_a875] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1976_c7_b851] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1983_c7_a875] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_return_output;

     -- t16_MUX[uxn_opcodes_h_l1976_c7_b851] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1976_c7_b851_cond <= VAR_t16_MUX_uxn_opcodes_h_l1976_c7_b851_cond;
     t16_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue;
     t16_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1976_c7_b851_return_output := t16_MUX_uxn_opcodes_h_l1976_c7_b851_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1983_c7_a875] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1976_c7_b851] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1976_c7_b851] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_return_output := result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1972_c7_5c34] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_a875_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1976_c7_b851_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1983_c7_a875_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_a875_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1976_c7_b851_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1976_c7_b851_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1976_c7_b851_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1976_c7_b851] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1976_c7_b851] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1972_c7_5c34] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output := result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1964_c2_c167] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1972_c7_5c34] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1972_c7_5c34] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output;

     -- t16_MUX[uxn_opcodes_h_l1972_c7_5c34] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1972_c7_5c34_cond <= VAR_t16_MUX_uxn_opcodes_h_l1972_c7_5c34_cond;
     t16_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue;
     t16_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output := t16_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1976_c7_b851] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1976_c7_b851_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1976_c7_b851_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1976_c7_b851_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1972_c7_5c34] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1964_c2_c167] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1972_c7_5c34] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1972_c7_5c34] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1964_c2_c167] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_return_output := result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_return_output;

     -- t16_MUX[uxn_opcodes_h_l1964_c2_c167] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1964_c2_c167_cond <= VAR_t16_MUX_uxn_opcodes_h_l1964_c2_c167_cond;
     t16_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue;
     t16_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1964_c2_c167_return_output := t16_MUX_uxn_opcodes_h_l1964_c2_c167_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1964_c2_c167] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_5c34_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l1964_c2_c167_return_output;
     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1964_c2_c167] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1964_c2_c167] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1964_c2_c167] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_return_output;

     -- Submodule level 5
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1989_l1960_DUPLICATE_9348 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1989_l1960_DUPLICATE_9348_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8152(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c2_c167_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c2_c167_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1964_c2_c167_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1964_c2_c167_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c2_c167_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c2_c167_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c2_c167_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1989_l1960_DUPLICATE_9348_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1989_l1960_DUPLICATE_9348_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
