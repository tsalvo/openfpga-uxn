-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 49
entity dei_0CLK_9bcaee2f is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_device_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dei_0CLK_9bcaee2f;
architecture arch of dei_0CLK_9bcaee2f is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal has_written_to_t : unsigned(0 downto 0) := to_unsigned(0, 1);
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal device_in_result : device_in_result_t := device_in_result_t_NULL;
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_has_written_to_t : unsigned(0 downto 0);
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_device_in_result : device_in_result_t;
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l403_c6_987e]
signal BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l419_c7_3235]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l403_c2_5333]
signal t8_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(7 downto 0);

-- device_in_result_MUX[uxn_opcodes_h_l403_c2_5333]
signal device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
signal device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_return_output : device_in_result_t;

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l403_c2_5333]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_return_output : signed(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l403_c2_5333]
signal result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l403_c2_5333]
signal result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l403_c2_5333]
signal result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(0 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l403_c2_5333]
signal result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l403_c2_5333]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l403_c2_5333]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l403_c2_5333]
signal result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l403_c2_5333]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(0 downto 0);

-- result_is_device_ram_write_MUX[uxn_opcodes_h_l403_c2_5333]
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l403_c2_5333]
signal result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(0 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l403_c2_5333]
signal has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l419_c11_01ff]
signal BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l422_c1_5d0f]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l419_c7_3235]
signal t8_MUX_uxn_opcodes_h_l419_c7_3235_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l419_c7_3235_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l419_c7_3235_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l419_c7_3235_return_output : unsigned(7 downto 0);

-- device_in_result_MUX[uxn_opcodes_h_l419_c7_3235]
signal device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_cond : unsigned(0 downto 0);
signal device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_iftrue : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_iffalse : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_return_output : device_in_result_t;

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l419_c7_3235]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l419_c7_3235]
signal result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l419_c7_3235]
signal result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l419_c7_3235]
signal result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_return_output : unsigned(0 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l419_c7_3235]
signal result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l419_c7_3235]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_return_output : unsigned(3 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l419_c7_3235]
signal has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l420_c30_7643]
signal sp_relative_shift_uxn_opcodes_h_l420_c30_7643_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l420_c30_7643_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l420_c30_7643_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l420_c30_7643_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l424_c9_74ec]
signal BIN_OP_EQ_uxn_opcodes_h_l424_c9_74ec_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l424_c9_74ec_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l424_c9_74ec_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l424_c9_6190]
signal MUX_uxn_opcodes_h_l424_c9_6190_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l424_c9_6190_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l424_c9_6190_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l424_c9_6190_return_output : unsigned(7 downto 0);

-- UNARY_OP_NOT[uxn_opcodes_h_l425_c8_edb7]
signal UNARY_OP_NOT_uxn_opcodes_h_l425_c8_edb7_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_uxn_opcodes_h_l425_c8_edb7_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l425_c1_e27e]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_return_output : unsigned(0 downto 0);

-- device_in_result_MUX[uxn_opcodes_h_l425_c3_a906]
signal device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_cond : unsigned(0 downto 0);
signal device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_iftrue : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_iffalse : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_return_output : device_in_result_t;

-- result_u8_value_MUX[uxn_opcodes_h_l425_c3_a906]
signal result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l425_c3_a906]
signal result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l425_c3_a906]
signal result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_return_output : unsigned(0 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l425_c3_a906]
signal result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l425_c3_a906]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_return_output : unsigned(3 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l425_c3_a906]
signal has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_return_output : unsigned(0 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_h_l426_c37_6593]
signal BIN_OP_MINUS_uxn_opcodes_h_l426_c37_6593_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l426_c37_6593_right : unsigned(1 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l426_c37_6593_return_output : unsigned(7 downto 0);

-- device_in[uxn_opcodes_h_l426_c23_f24d]
signal device_in_uxn_opcodes_h_l426_c23_f24d_CLOCK_ENABLE : unsigned(0 downto 0);
signal device_in_uxn_opcodes_h_l426_c23_f24d_device_address : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l426_c23_f24d_phase : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l426_c23_f24d_previous_device_ram_read : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l426_c23_f24d_return_output : device_in_result_t;

-- UNARY_OP_NOT[uxn_opcodes_h_l429_c9_72ee]
signal UNARY_OP_NOT_uxn_opcodes_h_l429_c9_72ee_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_uxn_opcodes_h_l429_c9_72ee_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l429_c4_d305]
signal result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l429_c4_d305]
signal result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l429_c4_d305]
signal result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l429_c4_d305]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_return_output : unsigned(3 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l429_c4_d305]
signal has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_return_output : unsigned(0 downto 0);

function CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6( ref_toks_0 : device_in_result_t;
 ref_toks_1 : unsigned) return device_in_result_t is
 
  variable base : device_in_result_t; 
  variable return_output : device_in_result_t;
begin
      base := ref_toks_0;
      base.is_dei_done := ref_toks_1;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_c644( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.device_ram_address := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;
      base.is_stack_index_flipped := ref_toks_7;
      base.u8_value := ref_toks_8;
      base.is_pc_updated := ref_toks_9;
      base.is_device_ram_write := ref_toks_10;
      base.is_vram_write := ref_toks_11;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e
BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_left,
BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_right,
BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_return_output);

-- t8_MUX_uxn_opcodes_h_l403_c2_5333
t8_MUX_uxn_opcodes_h_l403_c2_5333 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l403_c2_5333_cond,
t8_MUX_uxn_opcodes_h_l403_c2_5333_iftrue,
t8_MUX_uxn_opcodes_h_l403_c2_5333_iffalse,
t8_MUX_uxn_opcodes_h_l403_c2_5333_return_output);

-- device_in_result_MUX_uxn_opcodes_h_l403_c2_5333
device_in_result_MUX_uxn_opcodes_h_l403_c2_5333 : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_cond,
device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_iftrue,
device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_iffalse,
device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333
result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_cond,
result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_return_output);

-- result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_cond,
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_iftrue,
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_iffalse,
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_cond,
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff
BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_left,
BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_right,
BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_return_output);

-- t8_MUX_uxn_opcodes_h_l419_c7_3235
t8_MUX_uxn_opcodes_h_l419_c7_3235 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l419_c7_3235_cond,
t8_MUX_uxn_opcodes_h_l419_c7_3235_iftrue,
t8_MUX_uxn_opcodes_h_l419_c7_3235_iffalse,
t8_MUX_uxn_opcodes_h_l419_c7_3235_return_output);

-- device_in_result_MUX_uxn_opcodes_h_l419_c7_3235
device_in_result_MUX_uxn_opcodes_h_l419_c7_3235 : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_cond,
device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_iftrue,
device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_iffalse,
device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235
result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_cond,
result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_cond,
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_return_output);

-- sp_relative_shift_uxn_opcodes_h_l420_c30_7643
sp_relative_shift_uxn_opcodes_h_l420_c30_7643 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l420_c30_7643_ins,
sp_relative_shift_uxn_opcodes_h_l420_c30_7643_x,
sp_relative_shift_uxn_opcodes_h_l420_c30_7643_y,
sp_relative_shift_uxn_opcodes_h_l420_c30_7643_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l424_c9_74ec
BIN_OP_EQ_uxn_opcodes_h_l424_c9_74ec : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l424_c9_74ec_left,
BIN_OP_EQ_uxn_opcodes_h_l424_c9_74ec_right,
BIN_OP_EQ_uxn_opcodes_h_l424_c9_74ec_return_output);

-- MUX_uxn_opcodes_h_l424_c9_6190
MUX_uxn_opcodes_h_l424_c9_6190 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l424_c9_6190_cond,
MUX_uxn_opcodes_h_l424_c9_6190_iftrue,
MUX_uxn_opcodes_h_l424_c9_6190_iffalse,
MUX_uxn_opcodes_h_l424_c9_6190_return_output);

-- UNARY_OP_NOT_uxn_opcodes_h_l425_c8_edb7
UNARY_OP_NOT_uxn_opcodes_h_l425_c8_edb7 : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_uxn_opcodes_h_l425_c8_edb7_expr,
UNARY_OP_NOT_uxn_opcodes_h_l425_c8_edb7_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_return_output);

-- device_in_result_MUX_uxn_opcodes_h_l425_c3_a906
device_in_result_MUX_uxn_opcodes_h_l425_c3_a906 : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_cond,
device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_iftrue,
device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_iffalse,
device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906
result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_cond,
result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_cond,
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l426_c37_6593
BIN_OP_MINUS_uxn_opcodes_h_l426_c37_6593 : entity work.BIN_OP_MINUS_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l426_c37_6593_left,
BIN_OP_MINUS_uxn_opcodes_h_l426_c37_6593_right,
BIN_OP_MINUS_uxn_opcodes_h_l426_c37_6593_return_output);

-- device_in_uxn_opcodes_h_l426_c23_f24d
device_in_uxn_opcodes_h_l426_c23_f24d : entity work.device_in_0CLK_c6b159da port map (
clk,
device_in_uxn_opcodes_h_l426_c23_f24d_CLOCK_ENABLE,
device_in_uxn_opcodes_h_l426_c23_f24d_device_address,
device_in_uxn_opcodes_h_l426_c23_f24d_phase,
device_in_uxn_opcodes_h_l426_c23_f24d_previous_device_ram_read,
device_in_uxn_opcodes_h_l426_c23_f24d_return_output);

-- UNARY_OP_NOT_uxn_opcodes_h_l429_c9_72ee
UNARY_OP_NOT_uxn_opcodes_h_l429_c9_72ee : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_uxn_opcodes_h_l429_c9_72ee_expr,
UNARY_OP_NOT_uxn_opcodes_h_l429_c9_72ee_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305
result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_cond,
result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_cond,
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_device_ram_read,
 -- Registers
 has_written_to_t,
 t8,
 device_in_result,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_return_output,
 t8_MUX_uxn_opcodes_h_l403_c2_5333_return_output,
 device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_return_output,
 result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_return_output,
 t8_MUX_uxn_opcodes_h_l419_c7_3235_return_output,
 device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_return_output,
 sp_relative_shift_uxn_opcodes_h_l420_c30_7643_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l424_c9_74ec_return_output,
 MUX_uxn_opcodes_h_l424_c9_6190_return_output,
 UNARY_OP_NOT_uxn_opcodes_h_l425_c8_edb7_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_return_output,
 device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l426_c37_6593_return_output,
 device_in_uxn_opcodes_h_l426_c23_f24d_return_output,
 UNARY_OP_NOT_uxn_opcodes_h_l429_c9_72ee_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l419_c7_3235_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : device_in_result_t;
 variable VAR_device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6_uxn_opcodes_h_l403_c2_5333_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l408_c3_f682 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l414_c3_bd75 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l419_c7_3235_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l419_c7_3235_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l419_c7_3235_cond : unsigned(0 downto 0);
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_iftrue : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_iffalse : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l423_c3_cf80 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_cond : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_7643_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_7643_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_7643_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_7643_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l424_c9_6190_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_74ec_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_74ec_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_74ec_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l424_c9_6190_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l424_c9_6190_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l424_c9_6190_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d_uxn_opcodes_h_l425_c8_9390_return_output : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_edb7_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_edb7_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_iffalse : unsigned(0 downto 0);
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_iftrue : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_iffalse : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_cond : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_cond : unsigned(0 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_f24d_device_address : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_f24d_phase : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_f24d_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_6593_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_6593_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_6593_return_output : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_f24d_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_f24d_return_output : device_in_result_t;
 variable VAR_CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d_uxn_opcodes_h_l427_c32_1e19_return_output : unsigned(7 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_72ee_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_72ee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l431_c5_e71e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_cond : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d_uxn_opcodes_h_l432_c23_05f1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l425_l403_l419_DUPLICATE_c857_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l425_l403_l429_l419_DUPLICATE_652a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l425_l419_DUPLICATE_efe5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l425_l429_l419_DUPLICATE_4dd6_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l425_l429_l419_DUPLICATE_ce1f_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c644_uxn_opcodes_h_l441_l397_DUPLICATE_0906_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_has_written_to_t : unsigned(0 downto 0);
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_device_in_result : device_in_result_t;
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_has_written_to_t := has_written_to_t;
  REG_VAR_t8 := t8;
  REG_VAR_device_in_result := device_in_result;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_sp_relative_shift_uxn_opcodes_h_l423_c3_cf80 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_iffalse := VAR_result_sp_relative_shift_uxn_opcodes_h_l423_c3_cf80;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_iftrue := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_7643_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_iftrue := to_unsigned(1, 1);
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l414_c3_bd75 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l414_c3_bd75;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_right := to_unsigned(0, 1);
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_6593_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_iffalse := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_74ec_right := to_unsigned(2, 2);
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_7643_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l431_c5_e71e := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l431_c5_e71e;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l408_c3_f682 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l408_c3_f682;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_iftrue := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_right := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_device_ram_read := previous_device_ram_read;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_iffalse := VAR_CLOCK_ENABLE;
     VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_iftrue := device_in_result;
     VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_iffalse := device_in_result;
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_72ee_expr := has_written_to_t;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_iftrue := has_written_to_t;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_iftrue := has_written_to_t;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_iffalse := has_written_to_t;
     VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_7643_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_74ec_left := VAR_phase;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_6593_left := VAR_phase;
     VAR_device_in_uxn_opcodes_h_l426_c23_f24d_previous_device_ram_read := VAR_previous_device_ram_read;
     VAR_MUX_uxn_opcodes_h_l424_c9_6190_iftrue := VAR_previous_stack_read;
     VAR_MUX_uxn_opcodes_h_l424_c9_6190_iffalse := t8;
     VAR_t8_MUX_uxn_opcodes_h_l403_c2_5333_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l419_c7_3235_iftrue := t8;
     -- BIN_OP_MINUS[uxn_opcodes_h_l426_c37_6593] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l426_c37_6593_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_6593_left;
     BIN_OP_MINUS_uxn_opcodes_h_l426_c37_6593_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_6593_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_6593_return_output := BIN_OP_MINUS_uxn_opcodes_h_l426_c37_6593_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l403_c2_5333] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l403_c2_5333_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l425_l403_l429_l419_DUPLICATE_652a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l425_l403_l429_l419_DUPLICATE_652a_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l425_l419_DUPLICATE_efe5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l425_l419_DUPLICATE_efe5_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l425_l403_l419_DUPLICATE_c857 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l425_l403_l419_DUPLICATE_c857_return_output := result.device_ram_address;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l425_l429_l419_DUPLICATE_ce1f LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l425_l429_l419_DUPLICATE_ce1f_return_output := result.stack_address_sp_offset;

     -- device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6[uxn_opcodes_h_l403_c2_5333] LATENCY=0
     VAR_device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6_uxn_opcodes_h_l403_c2_5333_return_output := CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6(
     device_in_result,
     to_unsigned(0, 1));

     -- CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d[uxn_opcodes_h_l425_c8_9390] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d_uxn_opcodes_h_l425_c8_9390_return_output := device_in_result.is_dei_done;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l403_c2_5333] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l403_c2_5333_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l424_c9_74ec] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l424_c9_74ec_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_74ec_left;
     BIN_OP_EQ_uxn_opcodes_h_l424_c9_74ec_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_74ec_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_74ec_return_output := BIN_OP_EQ_uxn_opcodes_h_l424_c9_74ec_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l403_c2_5333] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l403_c2_5333_return_output := result.is_ram_write;

     -- result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d[uxn_opcodes_h_l403_c2_5333] LATENCY=0
     VAR_result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l403_c2_5333_return_output := result.is_device_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l419_c11_01ff] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_left;
     BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_return_output := BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_return_output;

     -- CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d[uxn_opcodes_h_l432_c23_05f1] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d_uxn_opcodes_h_l432_c23_05f1_return_output := device_in_result.dei_value;

     -- sp_relative_shift[uxn_opcodes_h_l420_c30_7643] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l420_c30_7643_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_7643_ins;
     sp_relative_shift_uxn_opcodes_h_l420_c30_7643_x <= VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_7643_x;
     sp_relative_shift_uxn_opcodes_h_l420_c30_7643_y <= VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_7643_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_7643_return_output := sp_relative_shift_uxn_opcodes_h_l420_c30_7643_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l425_l429_l419_DUPLICATE_4dd6 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l425_l429_l419_DUPLICATE_4dd6_return_output := result.is_opc_done;

     -- UNARY_OP_NOT[uxn_opcodes_h_l429_c9_72ee] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_uxn_opcodes_h_l429_c9_72ee_expr <= VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_72ee_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_72ee_return_output := UNARY_OP_NOT_uxn_opcodes_h_l429_c9_72ee_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l403_c2_5333] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l403_c2_5333_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l403_c6_987e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_left;
     BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_return_output := BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_return_output;

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l403_c2_5333_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_987e_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l419_c7_3235_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_01ff_return_output;
     VAR_MUX_uxn_opcodes_h_l424_c9_6190_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_74ec_return_output;
     VAR_device_in_uxn_opcodes_h_l426_c23_f24d_phase := VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_6593_return_output;
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_edb7_expr := VAR_CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d_uxn_opcodes_h_l425_c8_9390_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l425_l429_l419_DUPLICATE_4dd6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l425_l429_l419_DUPLICATE_4dd6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l425_l429_l419_DUPLICATE_4dd6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l425_l419_DUPLICATE_efe5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l425_l419_DUPLICATE_efe5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l425_l429_l419_DUPLICATE_ce1f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l425_l429_l419_DUPLICATE_ce1f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l425_l429_l419_DUPLICATE_ce1f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_iftrue := VAR_CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d_uxn_opcodes_h_l432_c23_05f1_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l425_l403_l419_DUPLICATE_c857_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l425_l403_l419_DUPLICATE_c857_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l425_l403_l419_DUPLICATE_c857_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l425_l403_l429_l419_DUPLICATE_652a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l425_l403_l429_l419_DUPLICATE_652a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l425_l403_l429_l419_DUPLICATE_652a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l425_l403_l429_l419_DUPLICATE_652a_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_72ee_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_72ee_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_72ee_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_72ee_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_72ee_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_iftrue := VAR_device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6_uxn_opcodes_h_l403_c2_5333_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_iffalse := VAR_result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l403_c2_5333_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l403_c2_5333_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l403_c2_5333_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l403_c2_5333_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l403_c2_5333_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_7643_return_output;
     -- result_is_ram_write_MUX[uxn_opcodes_h_l403_c2_5333] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output;

     -- MUX[uxn_opcodes_h_l424_c9_6190] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l424_c9_6190_cond <= VAR_MUX_uxn_opcodes_h_l424_c9_6190_cond;
     MUX_uxn_opcodes_h_l424_c9_6190_iftrue <= VAR_MUX_uxn_opcodes_h_l424_c9_6190_iftrue;
     MUX_uxn_opcodes_h_l424_c9_6190_iffalse <= VAR_MUX_uxn_opcodes_h_l424_c9_6190_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l424_c9_6190_return_output := MUX_uxn_opcodes_h_l424_c9_6190_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l403_c2_5333] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l429_c4_d305] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_return_output := has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l419_c7_3235] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l429_c4_d305] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_cond;
     result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_return_output := result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l429_c4_d305] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l429_c4_d305] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l403_c2_5333] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output;

     -- UNARY_OP_NOT[uxn_opcodes_h_l425_c8_edb7] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_uxn_opcodes_h_l425_c8_edb7_expr <= VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_edb7_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_edb7_return_output := UNARY_OP_NOT_uxn_opcodes_h_l425_c8_edb7_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l403_c2_5333] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_return_output;

     -- result_is_device_ram_write_MUX[uxn_opcodes_h_l403_c2_5333] LATENCY=0
     -- Inputs
     result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_cond <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_cond;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_iftrue <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_iftrue;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_iffalse <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_iffalse;
     -- Outputs
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output := result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l419_c7_3235] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l429_c4_d305] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_3235_return_output;
     VAR_device_in_uxn_opcodes_h_l426_c23_f24d_device_address := VAR_MUX_uxn_opcodes_h_l424_c9_6190_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l419_c7_3235_iffalse := VAR_MUX_uxn_opcodes_h_l424_c9_6190_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_edb7_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_edb7_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_edb7_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_edb7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_edb7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_edb7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_edb7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_edb7_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_iffalse := VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_d305_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_d305_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_d305_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_3235_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_d305_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_d305_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l422_c1_5d0f] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_return_output;

     -- t8_MUX[uxn_opcodes_h_l419_c7_3235] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l419_c7_3235_cond <= VAR_t8_MUX_uxn_opcodes_h_l419_c7_3235_cond;
     t8_MUX_uxn_opcodes_h_l419_c7_3235_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l419_c7_3235_iftrue;
     t8_MUX_uxn_opcodes_h_l419_c7_3235_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l419_c7_3235_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l419_c7_3235_return_output := t8_MUX_uxn_opcodes_h_l419_c7_3235_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l425_c3_a906] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_return_output := has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l425_c3_a906] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_cond;
     result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_return_output := result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l403_c2_5333] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l425_c3_a906] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l425_c3_a906] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l425_c3_a906] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_return_output;

     -- Submodule level 3
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_5d0f_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_iffalse := VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_a906_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_a906_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_a906_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_a906_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_a906_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l403_c2_5333_iffalse := VAR_t8_MUX_uxn_opcodes_h_l419_c7_3235_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l419_c7_3235] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l419_c7_3235] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l419_c7_3235] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_return_output := has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_return_output;

     -- t8_MUX[uxn_opcodes_h_l403_c2_5333] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l403_c2_5333_cond <= VAR_t8_MUX_uxn_opcodes_h_l403_c2_5333_cond;
     t8_MUX_uxn_opcodes_h_l403_c2_5333_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l403_c2_5333_iftrue;
     t8_MUX_uxn_opcodes_h_l403_c2_5333_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l403_c2_5333_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l403_c2_5333_return_output := t8_MUX_uxn_opcodes_h_l403_c2_5333_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l419_c7_3235] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l419_c7_3235] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_cond;
     result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_return_output := result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l425_c1_e27e] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_return_output;

     -- Submodule level 4
     VAR_device_in_uxn_opcodes_h_l426_c23_f24d_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_e27e_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_iffalse := VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_3235_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_3235_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_3235_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_3235_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_3235_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l403_c2_5333_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l403_c2_5333] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_cond;
     result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_return_output := result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l403_c2_5333] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l403_c2_5333] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_return_output;

     -- device_in[uxn_opcodes_h_l426_c23_f24d] LATENCY=0
     -- Clock enable
     device_in_uxn_opcodes_h_l426_c23_f24d_CLOCK_ENABLE <= VAR_device_in_uxn_opcodes_h_l426_c23_f24d_CLOCK_ENABLE;
     -- Inputs
     device_in_uxn_opcodes_h_l426_c23_f24d_device_address <= VAR_device_in_uxn_opcodes_h_l426_c23_f24d_device_address;
     device_in_uxn_opcodes_h_l426_c23_f24d_phase <= VAR_device_in_uxn_opcodes_h_l426_c23_f24d_phase;
     device_in_uxn_opcodes_h_l426_c23_f24d_previous_device_ram_read <= VAR_device_in_uxn_opcodes_h_l426_c23_f24d_previous_device_ram_read;
     -- Outputs
     VAR_device_in_uxn_opcodes_h_l426_c23_f24d_return_output := device_in_uxn_opcodes_h_l426_c23_f24d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l403_c2_5333] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l403_c2_5333] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_return_output := has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_return_output;

     -- Submodule level 5
     VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_iftrue := VAR_device_in_uxn_opcodes_h_l426_c23_f24d_return_output;
     REG_VAR_has_written_to_t := VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_5333_return_output;
     -- CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d[uxn_opcodes_h_l427_c32_1e19] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d_uxn_opcodes_h_l427_c32_1e19_return_output := VAR_device_in_uxn_opcodes_h_l426_c23_f24d_return_output.device_ram_address;

     -- device_in_result_MUX[uxn_opcodes_h_l425_c3_a906] LATENCY=0
     -- Inputs
     device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_cond <= VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_cond;
     device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_iftrue <= VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_iftrue;
     device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_iffalse <= VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_iffalse;
     -- Outputs
     VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_return_output := device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_return_output;

     -- Submodule level 6
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_iftrue := VAR_CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d_uxn_opcodes_h_l427_c32_1e19_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_iffalse := VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_a906_return_output;
     -- result_device_ram_address_MUX[uxn_opcodes_h_l425_c3_a906] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_return_output;

     -- device_in_result_MUX[uxn_opcodes_h_l419_c7_3235] LATENCY=0
     -- Inputs
     device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_cond <= VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_cond;
     device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_iftrue <= VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_iftrue;
     device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_iffalse <= VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_iffalse;
     -- Outputs
     VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_return_output := device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_return_output;

     -- Submodule level 7
     VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_iffalse := VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_3235_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_a906_return_output;
     -- result_device_ram_address_MUX[uxn_opcodes_h_l419_c7_3235] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_return_output;

     -- device_in_result_MUX[uxn_opcodes_h_l403_c2_5333] LATENCY=0
     -- Inputs
     device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_cond <= VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_cond;
     device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_iftrue <= VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_iftrue;
     device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_iffalse <= VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_iffalse;
     -- Outputs
     VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_return_output := device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_return_output;

     -- Submodule level 8
     REG_VAR_device_in_result := VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_5333_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_3235_return_output;
     -- result_device_ram_address_MUX[uxn_opcodes_h_l403_c2_5333] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_return_output;

     -- Submodule level 9
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c644_uxn_opcodes_h_l441_l397_DUPLICATE_0906 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c644_uxn_opcodes_h_l441_l397_DUPLICATE_0906_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c644(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_5333_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_5333_return_output,
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_5333_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_5333_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_5333_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_5333_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_5333_return_output,
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_5333_return_output);

     -- Submodule level 10
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c644_uxn_opcodes_h_l441_l397_DUPLICATE_0906_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c644_uxn_opcodes_h_l441_l397_DUPLICATE_0906_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_has_written_to_t <= REG_VAR_has_written_to_t;
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_device_in_result <= REG_VAR_device_in_result;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     has_written_to_t <= REG_COMB_has_written_to_t;
     t8 <= REG_COMB_t8;
     device_in_result <= REG_COMB_device_in_result;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
