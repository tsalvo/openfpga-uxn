-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity sth_0CLK_7883ef49 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sth_0CLK_7883ef49;
architecture arch of sth_0CLK_7883ef49 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2345_c6_71da]
signal BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2345_c2_600f]
signal result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2345_c2_600f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2345_c2_600f]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2345_c2_600f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2345_c2_600f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2345_c2_600f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2345_c2_600f]
signal t8_MUX_uxn_opcodes_h_l2345_c2_600f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2345_c2_600f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2352_c11_df93]
signal BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2352_c7_da96]
signal result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2352_c7_da96]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2352_c7_da96]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2352_c7_da96]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2352_c7_da96]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2352_c7_da96]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2352_c7_da96]
signal t8_MUX_uxn_opcodes_h_l2352_c7_da96_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2352_c7_da96_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2355_c11_201f]
signal BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2355_c7_88b1]
signal result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2355_c7_88b1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2355_c7_88b1]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2355_c7_88b1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2355_c7_88b1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2355_c7_88b1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2355_c7_88b1]
signal t8_MUX_uxn_opcodes_h_l2355_c7_88b1_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2358_c30_e277]
signal sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2360_c11_9a38]
signal BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2360_c7_6a1d]
signal result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2360_c7_6a1d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2360_c7_6a1d]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2360_c7_6a1d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2360_c7_6a1d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2360_c7_6a1d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2367_c11_3fd0]
signal BIN_OP_EQ_uxn_opcodes_h_l2367_c11_3fd0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2367_c11_3fd0_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2367_c11_3fd0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2367_c7_b9b7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2367_c7_b9b7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2367_c7_b9b7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2367_c7_b9b7]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_2b2f( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da
BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_left,
BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_right,
BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f
result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f
result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f
result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_return_output);

-- t8_MUX_uxn_opcodes_h_l2345_c2_600f
t8_MUX_uxn_opcodes_h_l2345_c2_600f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2345_c2_600f_cond,
t8_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue,
t8_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse,
t8_MUX_uxn_opcodes_h_l2345_c2_600f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93
BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_left,
BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_right,
BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96
result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_cond,
result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96
result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96
result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96
result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_return_output);

-- t8_MUX_uxn_opcodes_h_l2352_c7_da96
t8_MUX_uxn_opcodes_h_l2352_c7_da96 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2352_c7_da96_cond,
t8_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue,
t8_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse,
t8_MUX_uxn_opcodes_h_l2352_c7_da96_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f
BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_left,
BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_right,
BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1
result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_cond,
result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1
result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1
result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1
result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output);

-- t8_MUX_uxn_opcodes_h_l2355_c7_88b1
t8_MUX_uxn_opcodes_h_l2355_c7_88b1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2355_c7_88b1_cond,
t8_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue,
t8_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse,
t8_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2358_c30_e277
sp_relative_shift_uxn_opcodes_h_l2358_c30_e277 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_ins,
sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_x,
sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_y,
sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38
BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38_left,
BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38_right,
BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d
result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond,
result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d
result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d
result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d
result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2367_c11_3fd0
BIN_OP_EQ_uxn_opcodes_h_l2367_c11_3fd0 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2367_c11_3fd0_left,
BIN_OP_EQ_uxn_opcodes_h_l2367_c11_3fd0_right,
BIN_OP_EQ_uxn_opcodes_h_l2367_c11_3fd0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7
result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7
result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7
result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_return_output,
 t8_MUX_uxn_opcodes_h_l2345_c2_600f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_return_output,
 t8_MUX_uxn_opcodes_h_l2352_c7_da96_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output,
 t8_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output,
 sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2367_c11_3fd0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2349_c3_274f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2352_c7_da96_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2345_c2_600f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2345_c2_600f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2353_c3_b3af : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2352_c7_da96_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2355_c7_88b1_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2364_c3_d661 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2362_c3_d133 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2367_c11_3fd0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2367_c11_3fd0_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2367_c11_3fd0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2368_c3_14b6 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2360_l2352_l2355_l2345_DUPLICATE_2eff_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2352_l2367_l2355_l2345_DUPLICATE_1e57_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2352_l2367_l2355_l2345_DUPLICATE_50ed_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2352_l2367_l2345_DUPLICATE_e080_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2360_l2352_l2367_l2355_DUPLICATE_e3bf_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2360_l2355_DUPLICATE_8ca6_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_2b2f_uxn_opcodes_h_l2374_l2341_DUPLICATE_add0_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_y := resize(to_signed(-1, 2), 4);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2368_c3_14b6 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2368_c3_14b6;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2364_c3_d661 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2364_c3_d661;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2362_c3_d133 := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2362_c3_d133;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_right := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2349_c3_274f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2349_c3_274f;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2367_c11_3fd0_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2353_c3_b3af := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2353_c3_b3af;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2367_c11_3fd0_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2352_c11_df93] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_left;
     BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_return_output := BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2358_c30_e277] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_ins;
     sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_x;
     sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_return_output := sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2367_c11_3fd0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2367_c11_3fd0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2367_c11_3fd0_left;
     BIN_OP_EQ_uxn_opcodes_h_l2367_c11_3fd0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2367_c11_3fd0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2367_c11_3fd0_return_output := BIN_OP_EQ_uxn_opcodes_h_l2367_c11_3fd0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2355_c11_201f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2352_l2367_l2355_l2345_DUPLICATE_50ed LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2352_l2367_l2355_l2345_DUPLICATE_50ed_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l2360_c11_9a38] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38_left;
     BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38_return_output := BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2360_l2355_DUPLICATE_8ca6 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2360_l2355_DUPLICATE_8ca6_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2360_l2352_l2367_l2355_DUPLICATE_e3bf LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2360_l2352_l2367_l2355_DUPLICATE_e3bf_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2360_l2352_l2355_l2345_DUPLICATE_2eff LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2360_l2352_l2355_l2345_DUPLICATE_2eff_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2352_l2367_l2355_l2345_DUPLICATE_1e57 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2352_l2367_l2355_l2345_DUPLICATE_1e57_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2345_c6_71da] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_left;
     BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_return_output := BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2352_l2367_l2345_DUPLICATE_e080 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2352_l2367_l2345_DUPLICATE_e080_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2345_c2_600f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2345_c6_71da_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2352_c7_da96_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_df93_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2355_c7_88b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2355_c11_201f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2360_c11_9a38_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2367_c11_3fd0_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2367_c11_3fd0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2367_c11_3fd0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2367_c11_3fd0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2352_l2367_l2345_DUPLICATE_e080_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2352_l2367_l2345_DUPLICATE_e080_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2352_l2367_l2345_DUPLICATE_e080_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2360_l2352_l2367_l2355_DUPLICATE_e3bf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2360_l2352_l2367_l2355_DUPLICATE_e3bf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2360_l2352_l2367_l2355_DUPLICATE_e3bf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2360_l2352_l2367_l2355_DUPLICATE_e3bf_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2352_l2367_l2355_l2345_DUPLICATE_50ed_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2352_l2367_l2355_l2345_DUPLICATE_50ed_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2352_l2367_l2355_l2345_DUPLICATE_50ed_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2352_l2367_l2355_l2345_DUPLICATE_50ed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2352_l2367_l2355_l2345_DUPLICATE_1e57_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2352_l2367_l2355_l2345_DUPLICATE_1e57_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2352_l2367_l2355_l2345_DUPLICATE_1e57_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2352_l2367_l2355_l2345_DUPLICATE_1e57_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2360_l2355_DUPLICATE_8ca6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2360_l2355_DUPLICATE_8ca6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2360_l2352_l2355_l2345_DUPLICATE_2eff_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2360_l2352_l2355_l2345_DUPLICATE_2eff_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2360_l2352_l2355_l2345_DUPLICATE_2eff_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2360_l2352_l2355_l2345_DUPLICATE_2eff_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2358_c30_e277_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2367_c7_b9b7] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2367_c7_b9b7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2360_c7_6a1d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output := result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2360_c7_6a1d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2367_c7_b9b7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2367_c7_b9b7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output;

     -- t8_MUX[uxn_opcodes_h_l2355_c7_88b1] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2355_c7_88b1_cond <= VAR_t8_MUX_uxn_opcodes_h_l2355_c7_88b1_cond;
     t8_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue;
     t8_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output := t8_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2367_c7_b9b7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2360_c7_6a1d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2355_c7_88b1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2360_c7_6a1d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2360_c7_6a1d] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output;

     -- t8_MUX[uxn_opcodes_h_l2352_c7_da96] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2352_c7_da96_cond <= VAR_t8_MUX_uxn_opcodes_h_l2352_c7_da96_cond;
     t8_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue;
     t8_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2352_c7_da96_return_output := t8_MUX_uxn_opcodes_h_l2352_c7_da96_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2355_c7_88b1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output := result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2360_c7_6a1d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2360_c7_6a1d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2352_c7_da96_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2355_c7_88b1] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output;

     -- t8_MUX[uxn_opcodes_h_l2345_c2_600f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2345_c2_600f_cond <= VAR_t8_MUX_uxn_opcodes_h_l2345_c2_600f_cond;
     t8_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue;
     t8_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2345_c2_600f_return_output := t8_MUX_uxn_opcodes_h_l2345_c2_600f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2355_c7_88b1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2352_c7_da96] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2352_c7_da96] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_return_output := result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2355_c7_88b1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2355_c7_88b1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2355_c7_88b1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2352_c7_da96_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2352_c7_da96_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2345_c2_600f_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2345_c2_600f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2352_c7_da96] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2352_c7_da96] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2352_c7_da96] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2345_c2_600f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2352_c7_da96] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_da96_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2352_c7_da96_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_da96_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2352_c7_da96_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2345_c2_600f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2345_c2_600f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2345_c2_600f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2345_c2_600f] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_2b2f_uxn_opcodes_h_l2374_l2341_DUPLICATE_add0 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_2b2f_uxn_opcodes_h_l2374_l2341_DUPLICATE_add0_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_2b2f(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2345_c2_600f_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2345_c2_600f_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2345_c2_600f_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2345_c2_600f_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2345_c2_600f_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2345_c2_600f_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_2b2f_uxn_opcodes_h_l2374_l2341_DUPLICATE_add0_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_2b2f_uxn_opcodes_h_l2374_l2341_DUPLICATE_add0_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
