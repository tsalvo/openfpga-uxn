-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 52
entity mul_0CLK_f62d646e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end mul_0CLK_f62d646e;
architecture arch of mul_0CLK_f62d646e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2092_c6_134d]
signal BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2092_c1_9084]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2092_c2_268c]
signal n8_MUX_uxn_opcodes_h_l2092_c2_268c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2092_c2_268c_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2092_c2_268c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2092_c2_268c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2092_c2_268c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2092_c2_268c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2092_c2_268c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2092_c2_268c]
signal result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2092_c2_268c]
signal t8_MUX_uxn_opcodes_h_l2092_c2_268c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2092_c2_268c_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l2093_c3_8bae[uxn_opcodes_h_l2093_c3_8bae]
signal printf_uxn_opcodes_h_l2093_c3_8bae_uxn_opcodes_h_l2093_c3_8bae_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2097_c11_eb0a]
signal BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2097_c7_051f]
signal n8_MUX_uxn_opcodes_h_l2097_c7_051f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2097_c7_051f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2097_c7_051f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2097_c7_051f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2097_c7_051f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2097_c7_051f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2097_c7_051f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2097_c7_051f]
signal result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2097_c7_051f]
signal t8_MUX_uxn_opcodes_h_l2097_c7_051f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2097_c7_051f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2100_c11_c9f0]
signal BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2100_c7_fc9d]
signal n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2100_c7_fc9d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2100_c7_fc9d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2100_c7_fc9d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2100_c7_fc9d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2100_c7_fc9d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2100_c7_fc9d]
signal result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2100_c7_fc9d]
signal t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2104_c11_71ce]
signal BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2104_c7_29f2]
signal n8_MUX_uxn_opcodes_h_l2104_c7_29f2_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2104_c7_29f2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2104_c7_29f2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2104_c7_29f2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2104_c7_29f2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2104_c7_29f2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2104_c7_29f2]
signal result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2107_c11_0d94]
signal BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2107_c7_94d8]
signal n8_MUX_uxn_opcodes_h_l2107_c7_94d8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2107_c7_94d8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2107_c7_94d8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2107_c7_94d8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2107_c7_94d8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2107_c7_94d8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2107_c7_94d8]
signal result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2110_c30_b37a]
signal sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_return_output : signed(3 downto 0);

-- BIN_OP_INFERRED_MULT[uxn_opcodes_h_l2113_c21_373d]
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2113_c21_373d_left : unsigned(7 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2113_c21_373d_right : unsigned(7 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2113_c21_373d_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2115_c11_9682]
signal BIN_OP_EQ_uxn_opcodes_h_l2115_c11_9682_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2115_c11_9682_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2115_c11_9682_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2115_c7_f0a2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2115_c7_f0a2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2115_c7_f0a2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8cda( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d
BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_left,
BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_right,
BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_return_output);

-- n8_MUX_uxn_opcodes_h_l2092_c2_268c
n8_MUX_uxn_opcodes_h_l2092_c2_268c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2092_c2_268c_cond,
n8_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue,
n8_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse,
n8_MUX_uxn_opcodes_h_l2092_c2_268c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c
result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c
result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c
result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c
result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_return_output);

-- t8_MUX_uxn_opcodes_h_l2092_c2_268c
t8_MUX_uxn_opcodes_h_l2092_c2_268c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2092_c2_268c_cond,
t8_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue,
t8_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse,
t8_MUX_uxn_opcodes_h_l2092_c2_268c_return_output);

-- printf_uxn_opcodes_h_l2093_c3_8bae_uxn_opcodes_h_l2093_c3_8bae
printf_uxn_opcodes_h_l2093_c3_8bae_uxn_opcodes_h_l2093_c3_8bae : entity work.printf_uxn_opcodes_h_l2093_c3_8bae_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2093_c3_8bae_uxn_opcodes_h_l2093_c3_8bae_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a
BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_left,
BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_right,
BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_return_output);

-- n8_MUX_uxn_opcodes_h_l2097_c7_051f
n8_MUX_uxn_opcodes_h_l2097_c7_051f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2097_c7_051f_cond,
n8_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue,
n8_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse,
n8_MUX_uxn_opcodes_h_l2097_c7_051f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f
result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f
result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f
result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f
result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_return_output);

-- t8_MUX_uxn_opcodes_h_l2097_c7_051f
t8_MUX_uxn_opcodes_h_l2097_c7_051f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2097_c7_051f_cond,
t8_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue,
t8_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse,
t8_MUX_uxn_opcodes_h_l2097_c7_051f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0
BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_left,
BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_right,
BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_return_output);

-- n8_MUX_uxn_opcodes_h_l2100_c7_fc9d
n8_MUX_uxn_opcodes_h_l2100_c7_fc9d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond,
n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue,
n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse,
n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d
result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d
result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d
result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d
result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d
result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond,
result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output);

-- t8_MUX_uxn_opcodes_h_l2100_c7_fc9d
t8_MUX_uxn_opcodes_h_l2100_c7_fc9d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond,
t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue,
t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse,
t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce
BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_left,
BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_right,
BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_return_output);

-- n8_MUX_uxn_opcodes_h_l2104_c7_29f2
n8_MUX_uxn_opcodes_h_l2104_c7_29f2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2104_c7_29f2_cond,
n8_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue,
n8_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse,
n8_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2
result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2
result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2
result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2
result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2
result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_cond,
result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94
BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_left,
BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_right,
BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_return_output);

-- n8_MUX_uxn_opcodes_h_l2107_c7_94d8
n8_MUX_uxn_opcodes_h_l2107_c7_94d8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2107_c7_94d8_cond,
n8_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue,
n8_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse,
n8_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8
result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8
result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8
result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8
result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8
result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_cond,
result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a
sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_ins,
sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_x,
sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_y,
sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_return_output);

-- BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2113_c21_373d
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2113_c21_373d : entity work.BIN_OP_INFERRED_MULT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2113_c21_373d_left,
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2113_c21_373d_right,
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2113_c21_373d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2115_c11_9682
BIN_OP_EQ_uxn_opcodes_h_l2115_c11_9682 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2115_c11_9682_left,
BIN_OP_EQ_uxn_opcodes_h_l2115_c11_9682_right,
BIN_OP_EQ_uxn_opcodes_h_l2115_c11_9682_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2
result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2
result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2
result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_return_output,
 n8_MUX_uxn_opcodes_h_l2092_c2_268c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_return_output,
 t8_MUX_uxn_opcodes_h_l2092_c2_268c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_return_output,
 n8_MUX_uxn_opcodes_h_l2097_c7_051f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_return_output,
 t8_MUX_uxn_opcodes_h_l2097_c7_051f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_return_output,
 n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output,
 t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_return_output,
 n8_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_return_output,
 n8_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output,
 sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_return_output,
 BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2113_c21_373d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2115_c11_9682_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2097_c7_051f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2092_c2_268c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2092_c2_268c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2094_c3_ea3f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2097_c7_051f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2092_c2_268c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2092_c2_268c_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2093_c3_8bae_uxn_opcodes_h_l2093_c3_8bae_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2097_c7_051f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2098_c3_33ab : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2097_c7_051f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2102_c3_5fe5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2104_c7_29f2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2105_c3_797c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2107_c7_94d8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2112_c3_5ac4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2107_c7_94d8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_uxn_opcodes_h_l2113_c3_d02c : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2113_c21_373d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2113_c21_373d_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2113_c21_373d_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2115_c11_9682_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2115_c11_9682_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2115_c11_9682_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2107_DUPLICATE_e36e_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2115_DUPLICATE_1912_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2115_DUPLICATE_d31b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2107_DUPLICATE_eb7e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2115_l2107_DUPLICATE_8c0b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l2121_l2088_DUPLICATE_8578_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2098_c3_33ab := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2098_c3_33ab;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2112_c3_5ac4 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2112_c3_5ac4;
     VAR_sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2102_c3_5fe5 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2102_c3_5fe5;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2115_c11_9682_right := to_unsigned(5, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2094_c3_ea3f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2094_c3_ea3f;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2105_c3_797c := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2105_c3_797c;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_iffalse := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_right := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2115_c11_9682_left := VAR_phase;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2113_c21_373d_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2113_c21_373d_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2097_c11_eb0a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2107_c7_94d8] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2107_c7_94d8_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2107_DUPLICATE_e36e LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2107_DUPLICATE_e36e_return_output := result.sp_relative_shift;

     -- BIN_OP_INFERRED_MULT[uxn_opcodes_h_l2113_c21_373d] LATENCY=0
     -- Inputs
     BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2113_c21_373d_left <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2113_c21_373d_left;
     BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2113_c21_373d_right <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2113_c21_373d_right;
     -- Outputs
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2113_c21_373d_return_output := BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2113_c21_373d_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2107_DUPLICATE_eb7e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2107_DUPLICATE_eb7e_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2115_l2107_DUPLICATE_8c0b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2115_l2107_DUPLICATE_8c0b_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2115_c11_9682] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2115_c11_9682_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2115_c11_9682_left;
     BIN_OP_EQ_uxn_opcodes_h_l2115_c11_9682_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2115_c11_9682_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2115_c11_9682_return_output := BIN_OP_EQ_uxn_opcodes_h_l2115_c11_9682_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2100_c11_c9f0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_left;
     BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_return_output := BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2107_c11_0d94] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_left;
     BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_return_output := BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2110_c30_b37a] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_ins;
     sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_x;
     sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_return_output := sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2115_DUPLICATE_1912 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2115_DUPLICATE_1912_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2115_DUPLICATE_d31b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2115_DUPLICATE_d31b_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2092_c6_134d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_left;
     BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_return_output := BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2104_c11_71ce] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_left;
     BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_return_output := BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2092_c2_268c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2092_c2_268c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2092_c6_134d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2097_c7_051f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2097_c7_051f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_eb0a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2100_c11_c9f0_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2104_c7_29f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2104_c11_71ce_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2107_c7_94d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2107_c11_0d94_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2115_c11_9682_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2115_c11_9682_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2115_c11_9682_return_output;
     VAR_result_u8_value_uxn_opcodes_h_l2113_c3_d02c := resize(VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2113_c21_373d_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2107_DUPLICATE_e36e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2107_DUPLICATE_e36e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2107_DUPLICATE_e36e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2107_DUPLICATE_e36e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2107_DUPLICATE_e36e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2115_l2107_DUPLICATE_8c0b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2115_l2107_DUPLICATE_8c0b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2115_l2107_DUPLICATE_8c0b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2115_l2107_DUPLICATE_8c0b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2115_l2107_DUPLICATE_8c0b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2115_DUPLICATE_1912_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2115_DUPLICATE_1912_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2115_DUPLICATE_1912_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2115_DUPLICATE_1912_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2115_DUPLICATE_1912_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2115_DUPLICATE_d31b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2115_DUPLICATE_d31b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2115_DUPLICATE_d31b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2115_DUPLICATE_d31b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2115_DUPLICATE_d31b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2107_DUPLICATE_eb7e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2107_DUPLICATE_eb7e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2107_DUPLICATE_eb7e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2107_DUPLICATE_eb7e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2104_l2100_l2097_l2092_l2107_DUPLICATE_eb7e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2107_c7_94d8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2110_c30_b37a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue := VAR_result_u8_value_uxn_opcodes_h_l2113_c3_d02c;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2115_c7_f0a2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2107_c7_94d8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output;

     -- t8_MUX[uxn_opcodes_h_l2100_c7_fc9d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond <= VAR_t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond;
     t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue;
     t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output := t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2115_c7_f0a2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_return_output;

     -- n8_MUX[uxn_opcodes_h_l2107_c7_94d8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2107_c7_94d8_cond <= VAR_n8_MUX_uxn_opcodes_h_l2107_c7_94d8_cond;
     n8_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue;
     n8_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output := n8_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2115_c7_f0a2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2107_c7_94d8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2092_c1_9084] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2107_c7_94d8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output := result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l2093_c3_8bae_uxn_opcodes_h_l2093_c3_8bae_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2092_c1_9084_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2115_c7_f0a2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2115_c7_f0a2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2115_c7_f0a2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output;
     -- printf_uxn_opcodes_h_l2093_c3_8bae[uxn_opcodes_h_l2093_c3_8bae] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2093_c3_8bae_uxn_opcodes_h_l2093_c3_8bae_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2093_c3_8bae_uxn_opcodes_h_l2093_c3_8bae_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- t8_MUX[uxn_opcodes_h_l2097_c7_051f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2097_c7_051f_cond <= VAR_t8_MUX_uxn_opcodes_h_l2097_c7_051f_cond;
     t8_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue;
     t8_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2097_c7_051f_return_output := t8_MUX_uxn_opcodes_h_l2097_c7_051f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2104_c7_29f2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2107_c7_94d8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output;

     -- n8_MUX[uxn_opcodes_h_l2104_c7_29f2] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2104_c7_29f2_cond <= VAR_n8_MUX_uxn_opcodes_h_l2104_c7_29f2_cond;
     n8_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue;
     n8_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output := n8_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2107_c7_94d8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2104_c7_29f2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output := result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2107_c7_94d8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2104_c7_29f2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2107_c7_94d8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2097_c7_051f_return_output;
     -- n8_MUX[uxn_opcodes_h_l2100_c7_fc9d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond <= VAR_n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond;
     n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue;
     n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output := n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2104_c7_29f2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2100_c7_fc9d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output;

     -- t8_MUX[uxn_opcodes_h_l2092_c2_268c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2092_c2_268c_cond <= VAR_t8_MUX_uxn_opcodes_h_l2092_c2_268c_cond;
     t8_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue;
     t8_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2092_c2_268c_return_output := t8_MUX_uxn_opcodes_h_l2092_c2_268c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2104_c7_29f2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2100_c7_fc9d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output := result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2104_c7_29f2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2100_c7_fc9d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2104_c7_29f2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2092_c2_268c_return_output;
     -- n8_MUX[uxn_opcodes_h_l2097_c7_051f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2097_c7_051f_cond <= VAR_n8_MUX_uxn_opcodes_h_l2097_c7_051f_cond;
     n8_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue;
     n8_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2097_c7_051f_return_output := n8_MUX_uxn_opcodes_h_l2097_c7_051f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2100_c7_fc9d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2097_c7_051f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2100_c7_fc9d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2097_c7_051f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2100_c7_fc9d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2097_c7_051f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2097_c7_051f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2100_c7_fc9d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_051f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_051f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c7_051f_return_output;
     -- n8_MUX[uxn_opcodes_h_l2092_c2_268c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2092_c2_268c_cond <= VAR_n8_MUX_uxn_opcodes_h_l2092_c2_268c_cond;
     n8_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue;
     n8_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2092_c2_268c_return_output := n8_MUX_uxn_opcodes_h_l2092_c2_268c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2092_c2_268c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2097_c7_051f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2097_c7_051f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2092_c2_268c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2097_c7_051f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2092_c2_268c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2092_c2_268c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_051f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c7_051f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_051f_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2092_c2_268c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2092_c2_268c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2092_c2_268c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l2121_l2088_DUPLICATE_8578 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l2121_l2088_DUPLICATE_8578_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8cda(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2092_c2_268c_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2092_c2_268c_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2092_c2_268c_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2092_c2_268c_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2092_c2_268c_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2092_c2_268c_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l2121_l2088_DUPLICATE_8578_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l2121_l2088_DUPLICATE_8578_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
