-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 54
entity swp_0CLK_b288bfb7 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end swp_0CLK_b288bfb7;
architecture arch of swp_0CLK_b288bfb7 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2713_c6_66ae]
signal BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2713_c2_b8b8]
signal n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2713_c2_b8b8]
signal t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2713_c2_b8b8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2713_c2_b8b8]
signal result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2713_c2_b8b8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2713_c2_b8b8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2713_c2_b8b8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2713_c2_b8b8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2718_c11_bee5]
signal BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2718_c7_e4f9]
signal n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2718_c7_e4f9]
signal t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2718_c7_e4f9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2718_c7_e4f9]
signal result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2718_c7_e4f9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2718_c7_e4f9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2718_c7_e4f9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2718_c7_e4f9]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2721_c11_c3f2]
signal BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2721_c7_0b4a]
signal n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2721_c7_0b4a]
signal t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2721_c7_0b4a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2721_c7_0b4a]
signal result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2721_c7_0b4a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2721_c7_0b4a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2721_c7_0b4a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2721_c7_0b4a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2725_c11_d53e]
signal BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2725_c7_0dbb]
signal n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2725_c7_0dbb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2725_c7_0dbb]
signal result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2725_c7_0dbb]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2725_c7_0dbb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2725_c7_0dbb]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2725_c7_0dbb]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2728_c11_3586]
signal BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2728_c7_0a61]
signal n8_MUX_uxn_opcodes_h_l2728_c7_0a61_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2728_c7_0a61]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2728_c7_0a61]
signal result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2728_c7_0a61]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2728_c7_0a61]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2728_c7_0a61]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2728_c7_0a61]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2731_c30_a004]
signal sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2736_c11_d5ac]
signal BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2736_c7_7b86]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2736_c7_7b86]
signal result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2736_c7_7b86]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2736_c7_7b86]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2736_c7_7b86]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2741_c11_436d]
signal BIN_OP_EQ_uxn_opcodes_h_l2741_c11_436d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2741_c11_436d_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2741_c11_436d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2741_c7_d528]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2741_c7_d528]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_3345( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae
BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_left,
BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_right,
BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_return_output);

-- n8_MUX_uxn_opcodes_h_l2713_c2_b8b8
n8_MUX_uxn_opcodes_h_l2713_c2_b8b8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond,
n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue,
n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse,
n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output);

-- t8_MUX_uxn_opcodes_h_l2713_c2_b8b8
t8_MUX_uxn_opcodes_h_l2713_c2_b8b8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond,
t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue,
t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse,
t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8
result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond,
result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8
result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8
result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8
result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8
result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5
BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_left,
BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_right,
BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_return_output);

-- n8_MUX_uxn_opcodes_h_l2718_c7_e4f9
n8_MUX_uxn_opcodes_h_l2718_c7_e4f9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond,
n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue,
n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse,
n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output);

-- t8_MUX_uxn_opcodes_h_l2718_c7_e4f9
t8_MUX_uxn_opcodes_h_l2718_c7_e4f9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond,
t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue,
t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse,
t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9
result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond,
result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9
result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9
result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9
result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9
result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2
BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_left,
BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_right,
BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_return_output);

-- n8_MUX_uxn_opcodes_h_l2721_c7_0b4a
n8_MUX_uxn_opcodes_h_l2721_c7_0b4a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond,
n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue,
n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse,
n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output);

-- t8_MUX_uxn_opcodes_h_l2721_c7_0b4a
t8_MUX_uxn_opcodes_h_l2721_c7_0b4a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond,
t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue,
t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse,
t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a
result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond,
result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a
result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a
result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a
result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a
result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e
BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_left,
BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_right,
BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_return_output);

-- n8_MUX_uxn_opcodes_h_l2725_c7_0dbb
n8_MUX_uxn_opcodes_h_l2725_c7_0dbb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond,
n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue,
n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse,
n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb
result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond,
result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb
result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb
result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb
result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb
result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586
BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_left,
BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_right,
BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_return_output);

-- n8_MUX_uxn_opcodes_h_l2728_c7_0a61
n8_MUX_uxn_opcodes_h_l2728_c7_0a61 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2728_c7_0a61_cond,
n8_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue,
n8_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse,
n8_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61
result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_cond,
result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61
result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61
result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61
result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61
result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2731_c30_a004
sp_relative_shift_uxn_opcodes_h_l2731_c30_a004 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_ins,
sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_x,
sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_y,
sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac
BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac_left,
BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac_right,
BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86
result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_cond,
result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86
result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86
result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86
result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2741_c11_436d
BIN_OP_EQ_uxn_opcodes_h_l2741_c11_436d : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2741_c11_436d_left,
BIN_OP_EQ_uxn_opcodes_h_l2741_c11_436d_right,
BIN_OP_EQ_uxn_opcodes_h_l2741_c11_436d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528
result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528
result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_return_output,
 n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output,
 t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_return_output,
 n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output,
 t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_return_output,
 n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output,
 t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_return_output,
 n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_return_output,
 n8_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output,
 sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2741_c11_436d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2715_c3_f90a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2719_c3_be70 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2723_c3_24a7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2726_c3_fc79 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2728_c7_0a61_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2733_c3_cd93 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2738_c3_c4c4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2736_c7_7b86_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2741_c11_436d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2741_c11_436d_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2741_c11_436d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2736_DUPLICATE_f044_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2741_l2736_DUPLICATE_b6bb_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2728_DUPLICATE_ef88_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2736_DUPLICATE_493e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2741_l2736_l2728_DUPLICATE_6d3e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2746_l2709_DUPLICATE_9b3b_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2719_c3_be70 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2719_c3_be70;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2733_c3_cd93 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2733_c3_cd93;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2723_c3_24a7 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2723_c3_24a7;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2715_c3_f90a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2715_c3_f90a;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2741_c11_436d_right := to_unsigned(6, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac_right := to_unsigned(5, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2738_c3_c4c4 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2738_c3_c4c4;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2726_c3_fc79 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2726_c3_fc79;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2741_c11_436d_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2721_c11_c3f2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_left;
     BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_return_output := BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2728_DUPLICATE_ef88 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2728_DUPLICATE_ef88_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2725_c11_d53e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2736_c11_d5ac] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac_left;
     BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac_return_output := BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2728_c11_3586] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_left;
     BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_return_output := BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2741_c11_436d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2741_c11_436d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2741_c11_436d_left;
     BIN_OP_EQ_uxn_opcodes_h_l2741_c11_436d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2741_c11_436d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2741_c11_436d_return_output := BIN_OP_EQ_uxn_opcodes_h_l2741_c11_436d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2718_c11_bee5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_left;
     BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_return_output := BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2741_l2736_l2728_DUPLICATE_6d3e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2741_l2736_l2728_DUPLICATE_6d3e_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2736_DUPLICATE_493e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2736_DUPLICATE_493e_return_output := result.is_sp_shift;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2736_c7_7b86] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2736_c7_7b86_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2736_DUPLICATE_f044 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2736_DUPLICATE_f044_return_output := result.u8_value;

     -- sp_relative_shift[uxn_opcodes_h_l2731_c30_a004] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_ins;
     sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_x;
     sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_return_output := sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2741_l2736_DUPLICATE_b6bb LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2741_l2736_DUPLICATE_b6bb_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2713_c6_66ae] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_left;
     BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_return_output := BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2713_c6_66ae_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_bee5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2721_c11_c3f2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_d53e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2728_c7_0a61_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2728_c11_3586_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2736_c11_d5ac_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2741_c11_436d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2741_c11_436d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2728_DUPLICATE_ef88_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2728_DUPLICATE_ef88_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2728_DUPLICATE_ef88_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2728_DUPLICATE_ef88_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2728_DUPLICATE_ef88_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2741_l2736_l2728_DUPLICATE_6d3e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2741_l2736_l2728_DUPLICATE_6d3e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2741_l2736_l2728_DUPLICATE_6d3e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2741_l2736_l2728_DUPLICATE_6d3e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2741_l2736_l2728_DUPLICATE_6d3e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2741_l2736_l2728_DUPLICATE_6d3e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2736_DUPLICATE_493e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2736_DUPLICATE_493e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2736_DUPLICATE_493e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2736_DUPLICATE_493e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2736_DUPLICATE_493e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2741_l2736_DUPLICATE_b6bb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2741_l2736_DUPLICATE_b6bb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2741_l2736_DUPLICATE_b6bb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2741_l2736_DUPLICATE_b6bb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2741_l2736_DUPLICATE_b6bb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2741_l2736_DUPLICATE_b6bb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2736_DUPLICATE_f044_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2736_DUPLICATE_f044_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2736_DUPLICATE_f044_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2736_DUPLICATE_f044_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2725_l2721_l2718_l2713_l2736_DUPLICATE_f044_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2736_c7_7b86_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2731_c30_a004_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2736_c7_7b86] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2728_c7_0a61] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2736_c7_7b86] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output := result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2741_c7_d528] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2741_c7_d528] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_return_output;

     -- n8_MUX[uxn_opcodes_h_l2728_c7_0a61] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2728_c7_0a61_cond <= VAR_n8_MUX_uxn_opcodes_h_l2728_c7_0a61_cond;
     n8_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue;
     n8_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output := n8_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2736_c7_7b86] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output;

     -- t8_MUX[uxn_opcodes_h_l2721_c7_0b4a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond <= VAR_t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond;
     t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue;
     t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output := t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2741_c7_d528_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2741_c7_d528_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output;
     -- t8_MUX[uxn_opcodes_h_l2718_c7_e4f9] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond <= VAR_t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond;
     t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue;
     t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output := t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2736_c7_7b86] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2728_c7_0a61] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2725_c7_0dbb] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2736_c7_7b86] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2728_c7_0a61] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output;

     -- n8_MUX[uxn_opcodes_h_l2725_c7_0dbb] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond <= VAR_n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond;
     n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue;
     n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output := n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2728_c7_0a61] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output := result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2736_c7_7b86_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2725_c7_0dbb] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output := result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output;

     -- n8_MUX[uxn_opcodes_h_l2721_c7_0b4a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond <= VAR_n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond;
     n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue;
     n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output := n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2725_c7_0dbb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2728_c7_0a61] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2725_c7_0dbb] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2728_c7_0a61] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2721_c7_0b4a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output;

     -- t8_MUX[uxn_opcodes_h_l2713_c2_b8b8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond <= VAR_t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond;
     t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue;
     t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output := t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2728_c7_0a61_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output;
     -- n8_MUX[uxn_opcodes_h_l2718_c7_e4f9] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond <= VAR_n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond;
     n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue;
     n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output := n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2718_c7_e4f9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2721_c7_0b4a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2721_c7_0b4a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2725_c7_0dbb] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2725_c7_0dbb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2721_c7_0b4a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output := result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_0dbb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2721_c7_0b4a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2718_c7_e4f9] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2718_c7_e4f9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output;

     -- n8_MUX[uxn_opcodes_h_l2713_c2_b8b8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond <= VAR_n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond;
     n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue;
     n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output := n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2713_c2_b8b8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2721_c7_0b4a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2718_c7_e4f9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output := result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2721_c7_0b4a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2713_c2_b8b8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2713_c2_b8b8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2718_c7_e4f9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2713_c2_b8b8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output := result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2718_c7_e4f9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output;

     -- Submodule level 7
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e4f9_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2713_c2_b8b8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2713_c2_b8b8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output;

     -- Submodule level 8
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2746_l2709_DUPLICATE_9b3b LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2746_l2709_DUPLICATE_9b3b_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_3345(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2713_c2_b8b8_return_output);

     -- Submodule level 9
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2746_l2709_DUPLICATE_9b3b_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2746_l2709_DUPLICATE_9b3b_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
