-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity sta_0CLK_bce25fe8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sta_0CLK_bce25fe8;
architecture arch of sta_0CLK_bce25fe8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2299_c6_e7a0]
signal BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2299_c2_9f57]
signal result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2299_c2_9f57]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2299_c2_9f57]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2299_c2_9f57]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2299_c2_9f57]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2299_c2_9f57]
signal result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2299_c2_9f57]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2299_c2_9f57]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2299_c2_9f57]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2299_c2_9f57]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2299_c2_9f57]
signal t16_MUX_uxn_opcodes_h_l2299_c2_9f57_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(15 downto 0);

-- n8_MUX[uxn_opcodes_h_l2299_c2_9f57]
signal n8_MUX_uxn_opcodes_h_l2299_c2_9f57_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2312_c11_1428]
signal BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2312_c7_f9bd]
signal result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2312_c7_f9bd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output : unsigned(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2312_c7_f9bd]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2312_c7_f9bd]
signal result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2312_c7_f9bd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2312_c7_f9bd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2312_c7_f9bd]
signal t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output : unsigned(15 downto 0);

-- n8_MUX[uxn_opcodes_h_l2312_c7_f9bd]
signal n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2315_c11_7b57]
signal BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2315_c7_04a6]
signal result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2315_c7_04a6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output : unsigned(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2315_c7_04a6]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2315_c7_04a6]
signal result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2315_c7_04a6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2315_c7_04a6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2315_c7_04a6]
signal t16_MUX_uxn_opcodes_h_l2315_c7_04a6_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output : unsigned(15 downto 0);

-- n8_MUX[uxn_opcodes_h_l2315_c7_04a6]
signal n8_MUX_uxn_opcodes_h_l2315_c7_04a6_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output : unsigned(7 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l2317_c3_6213]
signal CONST_SL_8_uxn_opcodes_h_l2317_c3_6213_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l2317_c3_6213_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2320_c11_2a0c]
signal BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2320_c7_1532]
signal result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2320_c7_1532]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2320_c7_1532]
signal result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2320_c7_1532]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2320_c7_1532]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2320_c7_1532]
signal t16_MUX_uxn_opcodes_h_l2320_c7_1532_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2320_c7_1532_return_output : unsigned(15 downto 0);

-- n8_MUX[uxn_opcodes_h_l2320_c7_1532]
signal n8_MUX_uxn_opcodes_h_l2320_c7_1532_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2320_c7_1532_return_output : unsigned(7 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l2321_c3_efa5]
signal BIN_OP_OR_uxn_opcodes_h_l2321_c3_efa5_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2321_c3_efa5_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2321_c3_efa5_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2323_c11_a8e5]
signal BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2323_c7_60c9]
signal result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2323_c7_60c9]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2323_c7_60c9]
signal result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2323_c7_60c9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2323_c7_60c9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2323_c7_60c9]
signal n8_MUX_uxn_opcodes_h_l2323_c7_60c9_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2325_c30_7ae2]
signal sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_return_output : signed(3 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_2c6d( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : signed;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_vram_write := ref_toks_4;
      base.is_stack_index_flipped := ref_toks_5;
      base.u16_value := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.sp_relative_shift := ref_toks_9;
      base.is_opc_done := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0
BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_left,
BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_right,
BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57
result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_cond,
result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57
result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57
result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57
result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_cond,
result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57
result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57
result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57
result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57
result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output);

-- t16_MUX_uxn_opcodes_h_l2299_c2_9f57
t16_MUX_uxn_opcodes_h_l2299_c2_9f57 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2299_c2_9f57_cond,
t16_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue,
t16_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse,
t16_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output);

-- n8_MUX_uxn_opcodes_h_l2299_c2_9f57
n8_MUX_uxn_opcodes_h_l2299_c2_9f57 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2299_c2_9f57_cond,
n8_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue,
n8_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse,
n8_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428
BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_left,
BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_right,
BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd
result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond,
result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd
result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd
result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond,
result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd
result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd
result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output);

-- t16_MUX_uxn_opcodes_h_l2312_c7_f9bd
t16_MUX_uxn_opcodes_h_l2312_c7_f9bd : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond,
t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue,
t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse,
t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output);

-- n8_MUX_uxn_opcodes_h_l2312_c7_f9bd
n8_MUX_uxn_opcodes_h_l2312_c7_f9bd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond,
n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue,
n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse,
n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57
BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_left,
BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_right,
BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6
result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_cond,
result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6
result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6
result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_cond,
result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output);

-- t16_MUX_uxn_opcodes_h_l2315_c7_04a6
t16_MUX_uxn_opcodes_h_l2315_c7_04a6 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2315_c7_04a6_cond,
t16_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue,
t16_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse,
t16_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output);

-- n8_MUX_uxn_opcodes_h_l2315_c7_04a6
n8_MUX_uxn_opcodes_h_l2315_c7_04a6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2315_c7_04a6_cond,
n8_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue,
n8_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse,
n8_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output);

-- CONST_SL_8_uxn_opcodes_h_l2317_c3_6213
CONST_SL_8_uxn_opcodes_h_l2317_c3_6213 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l2317_c3_6213_x,
CONST_SL_8_uxn_opcodes_h_l2317_c3_6213_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c
BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_left,
BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_right,
BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532
result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_cond,
result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532
result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532
result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_cond,
result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532
result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532
result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_return_output);

-- t16_MUX_uxn_opcodes_h_l2320_c7_1532
t16_MUX_uxn_opcodes_h_l2320_c7_1532 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2320_c7_1532_cond,
t16_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue,
t16_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse,
t16_MUX_uxn_opcodes_h_l2320_c7_1532_return_output);

-- n8_MUX_uxn_opcodes_h_l2320_c7_1532
n8_MUX_uxn_opcodes_h_l2320_c7_1532 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2320_c7_1532_cond,
n8_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue,
n8_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse,
n8_MUX_uxn_opcodes_h_l2320_c7_1532_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l2321_c3_efa5
BIN_OP_OR_uxn_opcodes_h_l2321_c3_efa5 : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l2321_c3_efa5_left,
BIN_OP_OR_uxn_opcodes_h_l2321_c3_efa5_right,
BIN_OP_OR_uxn_opcodes_h_l2321_c3_efa5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5
BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5_left,
BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5_right,
BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9
result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_cond,
result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9
result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9
result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_cond,
result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9
result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9
result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output);

-- n8_MUX_uxn_opcodes_h_l2323_c7_60c9
n8_MUX_uxn_opcodes_h_l2323_c7_60c9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2323_c7_60c9_cond,
n8_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue,
n8_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse,
n8_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2
sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_ins,
sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_x,
sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_y,
sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output,
 t16_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output,
 n8_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output,
 t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output,
 n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output,
 t16_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output,
 n8_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output,
 CONST_SL_8_uxn_opcodes_h_l2317_c3_6213_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_return_output,
 t16_MUX_uxn_opcodes_h_l2320_c7_1532_return_output,
 n8_MUX_uxn_opcodes_h_l2320_c7_1532_return_output,
 BIN_OP_OR_uxn_opcodes_h_l2321_c3_efa5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output,
 n8_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output,
 sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2309_c3_1517 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2304_c3_e14a : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2299_c2_9f57_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2299_c2_9f57_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2313_c3_6395 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2318_c3_1da1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2315_c7_04a6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2320_c7_1532_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2315_c7_04a6_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2320_c7_1532_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2315_c7_04a6_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2317_c3_6213_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2317_c3_6213_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2320_c7_1532_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2320_c7_1532_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2321_c3_efa5_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2321_c3_efa5_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2321_c3_efa5_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2323_c7_60c9_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2315_l2312_l2299_l2323_l2320_DUPLICATE_03d3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2315_l2312_l2299_l2323_l2320_DUPLICATE_a12e_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2312_l2323_l2315_l2320_DUPLICATE_b4a2_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2312_l2323_l2315_l2320_DUPLICATE_fe03_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2312_l2323_l2315_l2320_DUPLICATE_03a8_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2316_l2321_DUPLICATE_6d80_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_2c6d_uxn_opcodes_h_l2294_l2332_DUPLICATE_6413_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2313_c3_6395 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2313_c3_6395;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2309_c3_1517 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2309_c3_1517;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2304_c3_e14a := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2304_c3_e14a;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2318_c3_1da1 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2318_c3_1da1;
     VAR_sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_y := resize(to_signed(-3, 3), 4);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_right := to_unsigned(3, 2);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2321_c3_efa5_left := t16;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse := t16;
     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2315_l2312_l2299_l2323_l2320_DUPLICATE_03d3 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2315_l2312_l2299_l2323_l2320_DUPLICATE_03d3_return_output := result.u8_value;

     -- sp_relative_shift[uxn_opcodes_h_l2325_c30_7ae2] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_ins;
     sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_x;
     sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_return_output := sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2299_c2_9f57] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2299_c2_9f57_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2315_l2312_l2299_l2323_l2320_DUPLICATE_a12e LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2315_l2312_l2299_l2323_l2320_DUPLICATE_a12e_return_output := result.u16_value;

     -- result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d[uxn_opcodes_h_l2299_c2_9f57] LATENCY=0
     VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2299_c2_9f57_return_output := result.is_stack_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2299_c2_9f57] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2299_c2_9f57_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2312_l2323_l2315_l2320_DUPLICATE_fe03 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2312_l2323_l2315_l2320_DUPLICATE_fe03_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2299_c6_e7a0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_left;
     BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_return_output := BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2312_l2323_l2315_l2320_DUPLICATE_03a8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2312_l2323_l2315_l2320_DUPLICATE_03a8_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2323_c11_a8e5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5_left;
     BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5_return_output := BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2299_c2_9f57] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2299_c2_9f57_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2312_l2323_l2315_l2320_DUPLICATE_b4a2 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2312_l2323_l2315_l2320_DUPLICATE_b4a2_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2315_c11_7b57] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_left;
     BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_return_output := BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2312_c11_1428] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_left;
     BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_return_output := BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2315_c7_04a6] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2315_c7_04a6_return_output := result.stack_address_sp_offset;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2316_l2321_DUPLICATE_6d80 LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2316_l2321_DUPLICATE_6d80_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l2320_c11_2a0c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l2299_c2_9f57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2299_c2_9f57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2299_c6_e7a0_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_1428_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2315_c7_04a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2315_c7_04a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_7b57_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2320_c7_1532_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2320_c7_1532_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_2a0c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2323_c7_60c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_a8e5_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2321_c3_efa5_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2316_l2321_DUPLICATE_6d80_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l2317_c3_6213_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2316_l2321_DUPLICATE_6d80_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2312_l2323_l2315_l2320_DUPLICATE_fe03_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2312_l2323_l2315_l2320_DUPLICATE_fe03_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2312_l2323_l2315_l2320_DUPLICATE_fe03_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2312_l2323_l2315_l2320_DUPLICATE_fe03_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2315_l2312_l2299_l2323_l2320_DUPLICATE_a12e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2315_l2312_l2299_l2323_l2320_DUPLICATE_a12e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2315_l2312_l2299_l2323_l2320_DUPLICATE_a12e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2315_l2312_l2299_l2323_l2320_DUPLICATE_a12e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2315_l2312_l2299_l2323_l2320_DUPLICATE_a12e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2312_l2323_l2315_l2320_DUPLICATE_03a8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2312_l2323_l2315_l2320_DUPLICATE_03a8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2312_l2323_l2315_l2320_DUPLICATE_03a8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2312_l2323_l2315_l2320_DUPLICATE_03a8_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2312_l2323_l2315_l2320_DUPLICATE_b4a2_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2312_l2323_l2315_l2320_DUPLICATE_b4a2_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2312_l2323_l2315_l2320_DUPLICATE_b4a2_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2312_l2323_l2315_l2320_DUPLICATE_b4a2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2315_l2312_l2299_l2323_l2320_DUPLICATE_03d3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2315_l2312_l2299_l2323_l2320_DUPLICATE_03d3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2315_l2312_l2299_l2323_l2320_DUPLICATE_03d3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2315_l2312_l2299_l2323_l2320_DUPLICATE_03d3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2315_l2312_l2299_l2323_l2320_DUPLICATE_03d3_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2299_c2_9f57_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2299_c2_9f57_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse := VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2299_c2_9f57_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2299_c2_9f57_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2315_c7_04a6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2325_c30_7ae2_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2323_c7_60c9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2299_c2_9f57] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l2321_c3_efa5] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l2321_c3_efa5_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l2321_c3_efa5_left;
     BIN_OP_OR_uxn_opcodes_h_l2321_c3_efa5_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l2321_c3_efa5_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l2321_c3_efa5_return_output := BIN_OP_OR_uxn_opcodes_h_l2321_c3_efa5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2299_c2_9f57] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2323_c7_60c9] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2323_c7_60c9] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output := result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2299_c2_9f57] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2315_c7_04a6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2323_c7_60c9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2299_c2_9f57] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2323_c7_60c9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output := result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output;

     -- n8_MUX[uxn_opcodes_h_l2323_c7_60c9] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2323_c7_60c9_cond <= VAR_n8_MUX_uxn_opcodes_h_l2323_c7_60c9_cond;
     n8_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2323_c7_60c9_iftrue;
     n8_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2323_c7_60c9_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output := n8_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l2317_c3_6213] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l2317_c3_6213_x <= VAR_CONST_SL_8_uxn_opcodes_h_l2317_c3_6213_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l2317_c3_6213_return_output := CONST_SL_8_uxn_opcodes_h_l2317_c3_6213_return_output;

     -- Submodule level 2
     VAR_t16_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l2321_c3_efa5_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l2317_c3_6213_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_60c9_return_output;
     -- t16_MUX[uxn_opcodes_h_l2320_c7_1532] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2320_c7_1532_cond <= VAR_t16_MUX_uxn_opcodes_h_l2320_c7_1532_cond;
     t16_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue;
     t16_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2320_c7_1532_return_output := t16_MUX_uxn_opcodes_h_l2320_c7_1532_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2320_c7_1532] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2320_c7_1532] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_return_output := result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_return_output;

     -- n8_MUX[uxn_opcodes_h_l2320_c7_1532] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2320_c7_1532_cond <= VAR_n8_MUX_uxn_opcodes_h_l2320_c7_1532_cond;
     n8_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue;
     n8_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2320_c7_1532_return_output := n8_MUX_uxn_opcodes_h_l2320_c7_1532_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2320_c7_1532] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_return_output := result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2320_c7_1532] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2312_c7_f9bd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2320_c7_1532] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2320_c7_1532_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_1532_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2320_c7_1532_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_1532_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2320_c7_1532_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_1532_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2320_c7_1532_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2315_c7_04a6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output;

     -- n8_MUX[uxn_opcodes_h_l2315_c7_04a6] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2315_c7_04a6_cond <= VAR_n8_MUX_uxn_opcodes_h_l2315_c7_04a6_cond;
     n8_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue;
     n8_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output := n8_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2315_c7_04a6] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2315_c7_04a6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output;

     -- t16_MUX[uxn_opcodes_h_l2315_c7_04a6] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2315_c7_04a6_cond <= VAR_t16_MUX_uxn_opcodes_h_l2315_c7_04a6_cond;
     t16_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue;
     t16_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output := t16_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2315_c7_04a6] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output := result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2315_c7_04a6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output := result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2299_c2_9f57] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2315_c7_04a6_return_output;
     -- n8_MUX[uxn_opcodes_h_l2312_c7_f9bd] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond <= VAR_n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond;
     n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue;
     n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output := n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2312_c7_f9bd] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output := result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2312_c7_f9bd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2312_c7_f9bd] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2312_c7_f9bd] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output := result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2312_c7_f9bd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output;

     -- t16_MUX[uxn_opcodes_h_l2312_c7_f9bd] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond <= VAR_t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_cond;
     t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_iftrue;
     t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output := t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2312_c7_f9bd_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2299_c2_9f57] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2299_c2_9f57] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2299_c2_9f57] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output := result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output;

     -- n8_MUX[uxn_opcodes_h_l2299_c2_9f57] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2299_c2_9f57_cond <= VAR_n8_MUX_uxn_opcodes_h_l2299_c2_9f57_cond;
     n8_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue;
     n8_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output := n8_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output;

     -- t16_MUX[uxn_opcodes_h_l2299_c2_9f57] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2299_c2_9f57_cond <= VAR_t16_MUX_uxn_opcodes_h_l2299_c2_9f57_cond;
     t16_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue;
     t16_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output := t16_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2299_c2_9f57] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2299_c2_9f57] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output := result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_2c6d_uxn_opcodes_h_l2294_l2332_DUPLICATE_6413 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_2c6d_uxn_opcodes_h_l2294_l2332_DUPLICATE_6413_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_2c6d(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2299_c2_9f57_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_2c6d_uxn_opcodes_h_l2294_l2332_DUPLICATE_6413_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_2c6d_uxn_opcodes_h_l2294_l2332_DUPLICATE_6413_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
