-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 55
entity ldr_0CLK_a6885b22 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldr_0CLK_a6885b22;
architecture arch of ldr_0CLK_a6885b22 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1694_c6_01d3]
signal BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1694_c1_96a6]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1694_c2_dea4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1694_c2_dea4]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1694_c2_dea4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1694_c2_dea4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1694_c2_dea4]
signal result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1694_c2_dea4]
signal result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1694_c2_dea4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output : signed(3 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1694_c2_dea4]
signal tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1694_c2_dea4]
signal t8_MUX_uxn_opcodes_h_l1694_c2_dea4_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1695_c3_380a[uxn_opcodes_h_l1695_c3_380a]
signal printf_uxn_opcodes_h_l1695_c3_380a_uxn_opcodes_h_l1695_c3_380a_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1699_c11_54c2]
signal BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1699_c7_1617]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1699_c7_1617]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1699_c7_1617]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1699_c7_1617]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1699_c7_1617]
signal result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1699_c7_1617]
signal result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1699_c7_1617]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_return_output : signed(3 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1699_c7_1617]
signal tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1699_c7_1617]
signal t8_MUX_uxn_opcodes_h_l1699_c7_1617_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1699_c7_1617_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1702_c11_6121]
signal BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1702_c7_d0f8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1702_c7_d0f8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1702_c7_d0f8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1702_c7_d0f8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1702_c7_d0f8]
signal result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1702_c7_d0f8]
signal result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1702_c7_d0f8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output : signed(3 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1702_c7_d0f8]
signal tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1702_c7_d0f8]
signal t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1705_c30_ada5]
signal sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_return_output : signed(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1706_c22_f27a]
signal BIN_OP_PLUS_uxn_opcodes_h_l1706_c22_f27a_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1706_c22_f27a_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1706_c22_f27a_return_output : signed(17 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1708_c11_372c]
signal BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1708_c7_5da0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1708_c7_5da0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1708_c7_5da0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1708_c7_5da0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1708_c7_5da0]
signal result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1708_c7_5da0]
signal result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1708_c7_5da0]
signal tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output : unsigned(7 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1710_c22_1d3a]
signal BIN_OP_PLUS_uxn_opcodes_h_l1710_c22_1d3a_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1710_c22_1d3a_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1710_c22_1d3a_return_output : signed(17 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1712_c11_35a4]
signal BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1712_c7_738e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1712_c7_738e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1712_c7_738e]
signal result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1712_c7_738e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1712_c7_738e]
signal tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1718_c11_86d2]
signal BIN_OP_EQ_uxn_opcodes_h_l1718_c11_86d2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1718_c11_86d2_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1718_c11_86d2_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1718_c7_f071]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1718_c7_f071]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_return_output : unsigned(0 downto 0);

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_284d( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.u16_value := ref_toks_5;
      base.u8_value := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3
BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_left,
BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_right,
BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4
result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4
result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4
result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4
result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_cond,
result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4
result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_cond,
result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4
result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4
tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_cond,
tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue,
tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse,
tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output);

-- t8_MUX_uxn_opcodes_h_l1694_c2_dea4
t8_MUX_uxn_opcodes_h_l1694_c2_dea4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1694_c2_dea4_cond,
t8_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue,
t8_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse,
t8_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output);

-- printf_uxn_opcodes_h_l1695_c3_380a_uxn_opcodes_h_l1695_c3_380a
printf_uxn_opcodes_h_l1695_c3_380a_uxn_opcodes_h_l1695_c3_380a : entity work.printf_uxn_opcodes_h_l1695_c3_380a_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1695_c3_380a_uxn_opcodes_h_l1695_c3_380a_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2
BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_left,
BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_right,
BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617
result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617
result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617
result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617
result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_cond,
result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617
result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_cond,
result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617
result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1699_c7_1617
tmp8_MUX_uxn_opcodes_h_l1699_c7_1617 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_cond,
tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue,
tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse,
tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_return_output);

-- t8_MUX_uxn_opcodes_h_l1699_c7_1617
t8_MUX_uxn_opcodes_h_l1699_c7_1617 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1699_c7_1617_cond,
t8_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue,
t8_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse,
t8_MUX_uxn_opcodes_h_l1699_c7_1617_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121
BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_left,
BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_right,
BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8
result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8
result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8
result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8
result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond,
result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8
result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond,
result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8
result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8
tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond,
tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue,
tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse,
tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output);

-- t8_MUX_uxn_opcodes_h_l1702_c7_d0f8
t8_MUX_uxn_opcodes_h_l1702_c7_d0f8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond,
t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue,
t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse,
t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5
sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_ins,
sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_x,
sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_y,
sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1706_c22_f27a
BIN_OP_PLUS_uxn_opcodes_h_l1706_c22_f27a : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1706_c22_f27a_left,
BIN_OP_PLUS_uxn_opcodes_h_l1706_c22_f27a_right,
BIN_OP_PLUS_uxn_opcodes_h_l1706_c22_f27a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c
BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_left,
BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_right,
BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0
result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0
result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0
result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0
result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_cond,
result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0
result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_cond,
result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0
tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_cond,
tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue,
tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse,
tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1710_c22_1d3a
BIN_OP_PLUS_uxn_opcodes_h_l1710_c22_1d3a : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1710_c22_1d3a_left,
BIN_OP_PLUS_uxn_opcodes_h_l1710_c22_1d3a_right,
BIN_OP_PLUS_uxn_opcodes_h_l1710_c22_1d3a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4
BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4_left,
BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4_right,
BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e
result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e
result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_cond,
result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e
result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1712_c7_738e
tmp8_MUX_uxn_opcodes_h_l1712_c7_738e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_cond,
tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue,
tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse,
tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1718_c11_86d2
BIN_OP_EQ_uxn_opcodes_h_l1718_c11_86d2 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1718_c11_86d2_left,
BIN_OP_EQ_uxn_opcodes_h_l1718_c11_86d2_right,
BIN_OP_EQ_uxn_opcodes_h_l1718_c11_86d2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071
result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071
result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output,
 tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output,
 t8_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_return_output,
 tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_return_output,
 t8_MUX_uxn_opcodes_h_l1699_c7_1617_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output,
 tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output,
 t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output,
 sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1706_c22_f27a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output,
 tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1710_c22_1d3a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_return_output,
 tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1718_c11_86d2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_iffalse : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1696_c3_75c1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1699_c7_1617_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1694_c2_dea4_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1695_c3_380a_uxn_opcodes_h_l1695_c3_380a_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1700_c3_e35a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1699_c7_1617_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l1706_c3_9350 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1706_c22_f27a_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l1706_c27_6a73_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1706_c22_f27a_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1706_c22_f27a_return_output : signed(17 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l1710_c3_3f3a : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1710_c22_1d3a_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l1710_c27_6324_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1710_c22_1d3a_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1710_c22_1d3a_return_output : signed(17 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1715_c3_e656 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_86d2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_86d2_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_86d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1694_l1708_l1699_DUPLICATE_486a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1708_l1702_l1699_l1694_l1718_DUPLICATE_d29f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1694_l1708_l1699_DUPLICATE_9c69_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1708_l1702_l1699_l1694_l1712_DUPLICATE_4cc3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1702_l1694_l1699_DUPLICATE_0905_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1708_l1702_l1699_l1718_l1712_DUPLICATE_b63d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1702_l1708_l1712_DUPLICATE_6a28_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_284d_uxn_opcodes_h_l1723_l1690_DUPLICATE_7d42_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1715_c3_e656 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1715_c3_e656;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1696_c3_75c1 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1696_c3_75c1;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_86d2_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1700_c3_e35a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1700_c3_e35a;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_iffalse := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_ins := VAR_ins;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1706_c22_f27a_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1710_c22_1d3a_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_86d2_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse := tmp8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1718_c11_86d2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1718_c11_86d2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_86d2_left;
     BIN_OP_EQ_uxn_opcodes_h_l1718_c11_86d2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_86d2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_86d2_return_output := BIN_OP_EQ_uxn_opcodes_h_l1718_c11_86d2_return_output;

     -- CAST_TO_int8_t[uxn_opcodes_h_l1710_c27_6324] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l1710_c27_6324_return_output := CAST_TO_int8_t_uint8_t(
     t8);

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1694_l1708_l1699_DUPLICATE_486a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1694_l1708_l1699_DUPLICATE_486a_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1694_l1708_l1699_DUPLICATE_9c69 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1694_l1708_l1699_DUPLICATE_9c69_return_output := result.u16_value;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1702_l1708_l1712_DUPLICATE_6a28 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1702_l1708_l1712_DUPLICATE_6a28_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1699_c11_54c2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_left;
     BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_return_output := BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1702_c11_6121] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_left;
     BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_return_output := BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1702_l1694_l1699_DUPLICATE_0905 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1702_l1694_l1699_DUPLICATE_0905_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1708_l1702_l1699_l1694_l1718_DUPLICATE_d29f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1708_l1702_l1699_l1694_l1718_DUPLICATE_d29f_return_output := result.is_stack_write;

     -- sp_relative_shift[uxn_opcodes_h_l1705_c30_ada5] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_ins;
     sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_x;
     sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_return_output := sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1708_l1702_l1699_l1694_l1712_DUPLICATE_4cc3 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1708_l1702_l1699_l1694_l1712_DUPLICATE_4cc3_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1712_c11_35a4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4_left;
     BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4_return_output := BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1694_c6_01d3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_left;
     BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_return_output := BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1708_c11_372c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_return_output;

     -- CAST_TO_int8_t[uxn_opcodes_h_l1706_c27_6a73] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l1706_c27_6a73_return_output := CAST_TO_int8_t_uint8_t(
     VAR_previous_stack_read);

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1708_l1702_l1699_l1718_l1712_DUPLICATE_b63d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1708_l1702_l1699_l1718_l1712_DUPLICATE_b63d_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1694_c2_dea4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c6_01d3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1699_c7_1617_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1699_c11_54c2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1702_c11_6121_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1708_c11_372c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1712_c11_35a4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_86d2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_86d2_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1706_c22_f27a_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l1706_c27_6a73_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1710_c22_1d3a_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l1710_c27_6324_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1702_l1694_l1699_DUPLICATE_0905_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1702_l1694_l1699_DUPLICATE_0905_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1702_l1694_l1699_DUPLICATE_0905_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1694_l1708_l1699_DUPLICATE_9c69_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1694_l1708_l1699_DUPLICATE_9c69_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1694_l1708_l1699_DUPLICATE_9c69_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1708_l1702_l1699_l1718_l1712_DUPLICATE_b63d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1708_l1702_l1699_l1718_l1712_DUPLICATE_b63d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1708_l1702_l1699_l1718_l1712_DUPLICATE_b63d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1708_l1702_l1699_l1718_l1712_DUPLICATE_b63d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1708_l1702_l1699_l1718_l1712_DUPLICATE_b63d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1694_l1708_l1699_DUPLICATE_486a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1694_l1708_l1699_DUPLICATE_486a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1694_l1708_l1699_DUPLICATE_486a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1708_l1702_l1699_l1694_l1718_DUPLICATE_d29f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1708_l1702_l1699_l1694_l1718_DUPLICATE_d29f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1708_l1702_l1699_l1694_l1718_DUPLICATE_d29f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1708_l1702_l1699_l1694_l1718_DUPLICATE_d29f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1708_l1702_l1699_l1694_l1718_DUPLICATE_d29f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1702_l1708_l1712_DUPLICATE_6a28_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1702_l1708_l1712_DUPLICATE_6a28_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1702_l1708_l1712_DUPLICATE_6a28_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1708_l1702_l1699_l1694_l1712_DUPLICATE_4cc3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1708_l1702_l1699_l1694_l1712_DUPLICATE_4cc3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1708_l1702_l1699_l1694_l1712_DUPLICATE_4cc3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1708_l1702_l1699_l1694_l1712_DUPLICATE_4cc3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1708_l1702_l1699_l1694_l1712_DUPLICATE_4cc3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1705_c30_ada5_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1712_c7_738e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_return_output := result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1702_c7_d0f8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1708_c7_5da0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output;

     -- t8_MUX[uxn_opcodes_h_l1702_c7_d0f8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond <= VAR_t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond;
     t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue;
     t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output := t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1710_c22_1d3a] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1710_c22_1d3a_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1710_c22_1d3a_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1710_c22_1d3a_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1710_c22_1d3a_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1710_c22_1d3a_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1710_c22_1d3a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1712_c7_738e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1712_c7_738e] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_cond;
     tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_return_output := tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1718_c7_f071] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1706_c22_f27a] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1706_c22_f27a_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1706_c22_f27a_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1706_c22_f27a_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1706_c22_f27a_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1706_c22_f27a_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1706_c22_f27a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1718_c7_f071] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1694_c1_96a6] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_return_output;

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l1706_c3_9350 := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1706_c22_f27a_return_output)),16);
     VAR_result_u16_value_uxn_opcodes_h_l1710_c3_3f3a := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1710_c22_1d3a_return_output)),16);
     VAR_printf_uxn_opcodes_h_l1695_c3_380a_uxn_opcodes_h_l1695_c3_380a_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1694_c1_96a6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_f071_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1718_c7_f071_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1712_c7_738e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1712_c7_738e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1712_c7_738e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue := VAR_result_u16_value_uxn_opcodes_h_l1706_c3_9350;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue := VAR_result_u16_value_uxn_opcodes_h_l1710_c3_3f3a;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1708_c7_5da0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output;

     -- t8_MUX[uxn_opcodes_h_l1699_c7_1617] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1699_c7_1617_cond <= VAR_t8_MUX_uxn_opcodes_h_l1699_c7_1617_cond;
     t8_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue;
     t8_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1699_c7_1617_return_output := t8_MUX_uxn_opcodes_h_l1699_c7_1617_return_output;

     -- printf_uxn_opcodes_h_l1695_c3_380a[uxn_opcodes_h_l1695_c3_380a] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1695_c3_380a_uxn_opcodes_h_l1695_c3_380a_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1695_c3_380a_uxn_opcodes_h_l1695_c3_380a_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_u8_value_MUX[uxn_opcodes_h_l1708_c7_5da0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output := result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1708_c7_5da0] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output := result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1702_c7_d0f8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1699_c7_1617] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1712_c7_738e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1712_c7_738e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1708_c7_5da0] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_cond;
     tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output := tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1712_c7_738e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1712_c7_738e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1699_c7_1617_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1699_c7_1617_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1708_c7_5da0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1702_c7_d0f8] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output := result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1699_c7_1617] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1702_c7_d0f8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output := result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output;

     -- t8_MUX[uxn_opcodes_h_l1694_c2_dea4] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1694_c2_dea4_cond <= VAR_t8_MUX_uxn_opcodes_h_l1694_c2_dea4_cond;
     t8_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue;
     t8_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output := t8_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1708_c7_5da0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1702_c7_d0f8] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond;
     tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output := tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1694_c2_dea4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1702_c7_d0f8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1699_c7_1617_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1708_c7_5da0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1702_c7_d0f8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1699_c7_1617] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_return_output := result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1702_c7_d0f8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1699_c7_1617] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1694_c2_dea4] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1699_c7_1617] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_return_output := result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1699_c7_1617] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_cond;
     tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_return_output := tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1702_c7_d0f8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1699_c7_1617_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1699_c7_1617_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1699_c7_1617_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1699_c7_1617_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l1694_c2_dea4] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output := result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1699_c7_1617] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1694_c2_dea4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output := result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1694_c2_dea4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1694_c2_dea4] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_cond;
     tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output := tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1699_c7_1617] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1699_c7_1617_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1699_c7_1617_return_output;
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1694_c2_dea4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1694_c2_dea4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_284d_uxn_opcodes_h_l1723_l1690_DUPLICATE_7d42 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_284d_uxn_opcodes_h_l1723_l1690_DUPLICATE_7d42_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_284d(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c2_dea4_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_284d_uxn_opcodes_h_l1723_l1690_DUPLICATE_7d42_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_284d_uxn_opcodes_h_l1723_l1690_DUPLICATE_7d42_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
