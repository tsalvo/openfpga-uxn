-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 50
entity ora_0CLK_fedec265 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ora_0CLK_fedec265;
architecture arch of ora_0CLK_fedec265 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1043_c6_d2c4]
signal BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1043_c2_5420]
signal n8_MUX_uxn_opcodes_h_l1043_c2_5420_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1043_c2_5420_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1043_c2_5420]
signal t8_MUX_uxn_opcodes_h_l1043_c2_5420_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1043_c2_5420_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1043_c2_5420]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1043_c2_5420]
signal result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1043_c2_5420]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1043_c2_5420]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1043_c2_5420]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1043_c2_5420]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1048_c11_2ad0]
signal BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1048_c7_d2df]
signal n8_MUX_uxn_opcodes_h_l1048_c7_d2df_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1048_c7_d2df]
signal t8_MUX_uxn_opcodes_h_l1048_c7_d2df_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1048_c7_d2df]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1048_c7_d2df]
signal result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1048_c7_d2df]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1048_c7_d2df]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1048_c7_d2df]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1048_c7_d2df]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1051_c11_45ed]
signal BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1051_c7_10a2]
signal n8_MUX_uxn_opcodes_h_l1051_c7_10a2_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1051_c7_10a2]
signal t8_MUX_uxn_opcodes_h_l1051_c7_10a2_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1051_c7_10a2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1051_c7_10a2]
signal result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1051_c7_10a2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1051_c7_10a2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1051_c7_10a2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1051_c7_10a2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1055_c11_26ac]
signal BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1055_c7_4200]
signal n8_MUX_uxn_opcodes_h_l1055_c7_4200_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1055_c7_4200_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1055_c7_4200]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1055_c7_4200]
signal result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1055_c7_4200]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1055_c7_4200]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1055_c7_4200]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1055_c7_4200]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1058_c11_61d1]
signal BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1058_c7_0cec]
signal n8_MUX_uxn_opcodes_h_l1058_c7_0cec_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1058_c7_0cec]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1058_c7_0cec]
signal result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1058_c7_0cec]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1058_c7_0cec]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1058_c7_0cec]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1058_c7_0cec]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1061_c30_2b95]
signal sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_return_output : signed(3 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l1064_c21_2884]
signal BIN_OP_OR_uxn_opcodes_h_l1064_c21_2884_left : unsigned(7 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l1064_c21_2884_right : unsigned(7 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l1064_c21_2884_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1066_c11_17ea]
signal BIN_OP_EQ_uxn_opcodes_h_l1066_c11_17ea_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1066_c11_17ea_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1066_c11_17ea_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1066_c7_02ee]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1066_c7_02ee]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1066_c7_02ee]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_3345( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4
BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_left,
BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_right,
BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_return_output);

-- n8_MUX_uxn_opcodes_h_l1043_c2_5420
n8_MUX_uxn_opcodes_h_l1043_c2_5420 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1043_c2_5420_cond,
n8_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue,
n8_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse,
n8_MUX_uxn_opcodes_h_l1043_c2_5420_return_output);

-- t8_MUX_uxn_opcodes_h_l1043_c2_5420
t8_MUX_uxn_opcodes_h_l1043_c2_5420 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1043_c2_5420_cond,
t8_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue,
t8_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse,
t8_MUX_uxn_opcodes_h_l1043_c2_5420_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420
result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_cond,
result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420
result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420
result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420
result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420
result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0
BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_left,
BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_right,
BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_return_output);

-- n8_MUX_uxn_opcodes_h_l1048_c7_d2df
n8_MUX_uxn_opcodes_h_l1048_c7_d2df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1048_c7_d2df_cond,
n8_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue,
n8_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse,
n8_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output);

-- t8_MUX_uxn_opcodes_h_l1048_c7_d2df
t8_MUX_uxn_opcodes_h_l1048_c7_d2df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1048_c7_d2df_cond,
t8_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue,
t8_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse,
t8_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df
result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_cond,
result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df
result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df
result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df
result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df
result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed
BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_left,
BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_right,
BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_return_output);

-- n8_MUX_uxn_opcodes_h_l1051_c7_10a2
n8_MUX_uxn_opcodes_h_l1051_c7_10a2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1051_c7_10a2_cond,
n8_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue,
n8_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse,
n8_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output);

-- t8_MUX_uxn_opcodes_h_l1051_c7_10a2
t8_MUX_uxn_opcodes_h_l1051_c7_10a2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1051_c7_10a2_cond,
t8_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue,
t8_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse,
t8_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2
result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_cond,
result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2
result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2
result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2
result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2
result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac
BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_left,
BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_right,
BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_return_output);

-- n8_MUX_uxn_opcodes_h_l1055_c7_4200
n8_MUX_uxn_opcodes_h_l1055_c7_4200 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1055_c7_4200_cond,
n8_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue,
n8_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse,
n8_MUX_uxn_opcodes_h_l1055_c7_4200_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200
result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_cond,
result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200
result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200
result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200
result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200
result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1
BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_left,
BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_right,
BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_return_output);

-- n8_MUX_uxn_opcodes_h_l1058_c7_0cec
n8_MUX_uxn_opcodes_h_l1058_c7_0cec : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1058_c7_0cec_cond,
n8_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue,
n8_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse,
n8_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec
result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_cond,
result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec
result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec
result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec
result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec
result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95
sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_ins,
sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_x,
sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_y,
sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l1064_c21_2884
BIN_OP_OR_uxn_opcodes_h_l1064_c21_2884 : entity work.BIN_OP_OR_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l1064_c21_2884_left,
BIN_OP_OR_uxn_opcodes_h_l1064_c21_2884_right,
BIN_OP_OR_uxn_opcodes_h_l1064_c21_2884_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1066_c11_17ea
BIN_OP_EQ_uxn_opcodes_h_l1066_c11_17ea : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1066_c11_17ea_left,
BIN_OP_EQ_uxn_opcodes_h_l1066_c11_17ea_right,
BIN_OP_EQ_uxn_opcodes_h_l1066_c11_17ea_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee
result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee
result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee
result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_return_output,
 n8_MUX_uxn_opcodes_h_l1043_c2_5420_return_output,
 t8_MUX_uxn_opcodes_h_l1043_c2_5420_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_return_output,
 n8_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output,
 t8_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_return_output,
 n8_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output,
 t8_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_return_output,
 n8_MUX_uxn_opcodes_h_l1055_c7_4200_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_return_output,
 n8_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output,
 sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_return_output,
 BIN_OP_OR_uxn_opcodes_h_l1064_c21_2884_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1066_c11_17ea_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1043_c2_5420_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1043_c2_5420_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1043_c2_5420_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1043_c2_5420_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1045_c3_6004 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1048_c7_d2df_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1048_c7_d2df_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1049_c3_8b93 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1055_c7_4200_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1051_c7_10a2_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1051_c7_10a2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1053_c3_5ecf : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1055_c7_4200_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1056_c3_da25 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1058_c7_0cec_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1063_c3_921b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1058_c7_0cec_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1064_c21_2884_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1064_c21_2884_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1064_c21_2884_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1066_c11_17ea_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1066_c11_17ea_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1066_c11_17ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1058_DUPLICATE_4d53_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1066_DUPLICATE_8c90_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1058_DUPLICATE_655d_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1066_DUPLICATE_2153_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1066_l1058_DUPLICATE_0339_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1072_l1039_DUPLICATE_bd98_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1056_c3_da25 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1056_c3_da25;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1066_c11_17ea_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1063_c3_921b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1063_c3_921b;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1053_c3_5ecf := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1053_c3_5ecf;
     VAR_sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1049_c3_8b93 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1049_c3_8b93;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1045_c3_6004 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1045_c3_6004;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1066_c11_17ea_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l1064_c21_2884_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_OR_uxn_opcodes_h_l1064_c21_2884_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse := t8;
     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1058_c7_0cec] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1058_c7_0cec_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1066_DUPLICATE_8c90 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1066_DUPLICATE_8c90_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1066_c11_17ea] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1066_c11_17ea_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1066_c11_17ea_left;
     BIN_OP_EQ_uxn_opcodes_h_l1066_c11_17ea_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1066_c11_17ea_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1066_c11_17ea_return_output := BIN_OP_EQ_uxn_opcodes_h_l1066_c11_17ea_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1058_c11_61d1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_left;
     BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_return_output := BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1043_c6_d2c4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_left;
     BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_return_output := BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1061_c30_2b95] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_ins;
     sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_x;
     sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_return_output := sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1055_c11_26ac] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_left;
     BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_return_output := BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1058_DUPLICATE_655d LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1058_DUPLICATE_655d_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1058_DUPLICATE_4d53 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1058_DUPLICATE_4d53_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1066_DUPLICATE_2153 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1066_DUPLICATE_2153_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1066_l1058_DUPLICATE_0339 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1066_l1058_DUPLICATE_0339_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1048_c11_2ad0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_left;
     BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_return_output := BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1051_c11_45ed] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_left;
     BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_return_output := BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l1064_c21_2884] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l1064_c21_2884_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l1064_c21_2884_left;
     BIN_OP_OR_uxn_opcodes_h_l1064_c21_2884_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l1064_c21_2884_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l1064_c21_2884_return_output := BIN_OP_OR_uxn_opcodes_h_l1064_c21_2884_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1043_c2_5420_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1043_c2_5420_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c6_d2c4_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1048_c7_d2df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1048_c7_d2df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1048_c11_2ad0_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1051_c7_10a2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1051_c7_10a2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1051_c11_45ed_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1055_c7_4200_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1055_c11_26ac_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1058_c7_0cec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1058_c11_61d1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1066_c11_17ea_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1066_c11_17ea_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1066_c11_17ea_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l1064_c21_2884_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1058_DUPLICATE_655d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1058_DUPLICATE_655d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1058_DUPLICATE_655d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1058_DUPLICATE_655d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1058_DUPLICATE_655d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1066_l1058_DUPLICATE_0339_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1066_l1058_DUPLICATE_0339_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1066_l1058_DUPLICATE_0339_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1066_l1058_DUPLICATE_0339_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1066_l1058_DUPLICATE_0339_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1066_DUPLICATE_2153_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1066_DUPLICATE_2153_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1066_DUPLICATE_2153_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1066_DUPLICATE_2153_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1066_DUPLICATE_2153_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1066_DUPLICATE_8c90_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1066_DUPLICATE_8c90_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1066_DUPLICATE_8c90_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1066_DUPLICATE_8c90_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1066_DUPLICATE_8c90_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1058_DUPLICATE_4d53_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1058_DUPLICATE_4d53_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1058_DUPLICATE_4d53_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1058_DUPLICATE_4d53_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1055_l1051_l1048_l1043_l1058_DUPLICATE_4d53_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1058_c7_0cec_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1061_c30_2b95_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1058_c7_0cec] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output := result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1058_c7_0cec] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output;

     -- n8_MUX[uxn_opcodes_h_l1058_c7_0cec] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1058_c7_0cec_cond <= VAR_n8_MUX_uxn_opcodes_h_l1058_c7_0cec_cond;
     n8_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue;
     n8_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output := n8_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1066_c7_02ee] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_return_output;

     -- t8_MUX[uxn_opcodes_h_l1051_c7_10a2] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1051_c7_10a2_cond <= VAR_t8_MUX_uxn_opcodes_h_l1051_c7_10a2_cond;
     t8_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue;
     t8_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output := t8_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1066_c7_02ee] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1058_c7_0cec] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1066_c7_02ee] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1066_c7_02ee_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1066_c7_02ee_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1066_c7_02ee_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1058_c7_0cec] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1058_c7_0cec] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1055_c7_4200] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_return_output;

     -- n8_MUX[uxn_opcodes_h_l1055_c7_4200] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1055_c7_4200_cond <= VAR_n8_MUX_uxn_opcodes_h_l1055_c7_4200_cond;
     n8_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue;
     n8_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1055_c7_4200_return_output := n8_MUX_uxn_opcodes_h_l1055_c7_4200_return_output;

     -- t8_MUX[uxn_opcodes_h_l1048_c7_d2df] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1048_c7_d2df_cond <= VAR_t8_MUX_uxn_opcodes_h_l1048_c7_d2df_cond;
     t8_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue;
     t8_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output := t8_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1055_c7_4200] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_return_output := result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1055_c7_4200] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1058_c7_0cec] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1055_c7_4200_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1058_c7_0cec_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1055_c7_4200_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1055_c7_4200_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1055_c7_4200_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1055_c7_4200] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1051_c7_10a2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output := result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1055_c7_4200] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_return_output;

     -- t8_MUX[uxn_opcodes_h_l1043_c2_5420] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1043_c2_5420_cond <= VAR_t8_MUX_uxn_opcodes_h_l1043_c2_5420_cond;
     t8_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue;
     t8_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1043_c2_5420_return_output := t8_MUX_uxn_opcodes_h_l1043_c2_5420_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1051_c7_10a2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1055_c7_4200] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1051_c7_10a2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output;

     -- n8_MUX[uxn_opcodes_h_l1051_c7_10a2] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1051_c7_10a2_cond <= VAR_n8_MUX_uxn_opcodes_h_l1051_c7_10a2_cond;
     n8_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue;
     n8_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output := n8_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1055_c7_4200_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1055_c7_4200_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1055_c7_4200_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1043_c2_5420_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1048_c7_d2df] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1051_c7_10a2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1051_c7_10a2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1051_c7_10a2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1048_c7_d2df] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output;

     -- n8_MUX[uxn_opcodes_h_l1048_c7_d2df] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1048_c7_d2df_cond <= VAR_n8_MUX_uxn_opcodes_h_l1048_c7_d2df_cond;
     n8_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue;
     n8_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output := n8_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1048_c7_d2df] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output := result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1051_c7_10a2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1043_c2_5420] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_return_output;

     -- n8_MUX[uxn_opcodes_h_l1043_c2_5420] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1043_c2_5420_cond <= VAR_n8_MUX_uxn_opcodes_h_l1043_c2_5420_cond;
     n8_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue;
     n8_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1043_c2_5420_return_output := n8_MUX_uxn_opcodes_h_l1043_c2_5420_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1048_c7_d2df] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1048_c7_d2df] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1043_c2_5420] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_return_output := result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1048_c7_d2df] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1043_c2_5420] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1043_c2_5420_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1048_c7_d2df_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1043_c2_5420] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1043_c2_5420] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1043_c2_5420] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1072_l1039_DUPLICATE_bd98 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1072_l1039_DUPLICATE_bd98_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_3345(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c2_5420_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c2_5420_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c2_5420_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c2_5420_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c2_5420_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c2_5420_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1072_l1039_DUPLICATE_bd98_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1072_l1039_DUPLICATE_bd98_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
