-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 46
entity ldz_0CLK_fd0ee55b is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldz_0CLK_fd0ee55b;
architecture arch of ldz_0CLK_fd0ee55b is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1409_c6_4d0f]
signal BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1409_c2_b22e]
signal tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1409_c2_b22e]
signal result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1409_c2_b22e]
signal result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1409_c2_b22e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1409_c2_b22e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1409_c2_b22e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1409_c2_b22e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1409_c2_b22e]
signal t8_MUX_uxn_opcodes_h_l1409_c2_b22e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1416_c11_2f58]
signal BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1416_c7_b689]
signal tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1416_c7_b689]
signal result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1416_c7_b689]
signal result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1416_c7_b689]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1416_c7_b689]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1416_c7_b689]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1416_c7_b689]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1416_c7_b689]
signal t8_MUX_uxn_opcodes_h_l1416_c7_b689_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1416_c7_b689_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1419_c11_a6bb]
signal BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1419_c7_fa4b]
signal tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1419_c7_fa4b]
signal result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1419_c7_fa4b]
signal result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1419_c7_fa4b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1419_c7_fa4b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1419_c7_fa4b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1419_c7_fa4b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1419_c7_fa4b]
signal t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1422_c30_c99b]
signal sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1425_c11_72a3]
signal BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1425_c7_7691]
signal tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1425_c7_7691]
signal result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1425_c7_7691]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1425_c7_7691]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1425_c7_7691]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1425_c7_7691]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1428_c11_ba0b]
signal BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1428_c7_ad75]
signal tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1428_c7_ad75]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1428_c7_ad75]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1428_c7_ad75]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1428_c7_ad75]
signal result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1434_c11_6cab]
signal BIN_OP_EQ_uxn_opcodes_h_l1434_c11_6cab_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1434_c11_6cab_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1434_c11_6cab_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1434_c7_9420]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1434_c7_9420]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_return_output : unsigned(0 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_e78e( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u16_value := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f
BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_left,
BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_right,
BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e
tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_cond,
tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue,
tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse,
tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e
result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_cond,
result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e
result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_cond,
result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e
result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e
result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e
result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output);

-- t8_MUX_uxn_opcodes_h_l1409_c2_b22e
t8_MUX_uxn_opcodes_h_l1409_c2_b22e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1409_c2_b22e_cond,
t8_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue,
t8_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse,
t8_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58
BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_left,
BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_right,
BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1416_c7_b689
tmp8_MUX_uxn_opcodes_h_l1416_c7_b689 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_cond,
tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue,
tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse,
tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689
result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_cond,
result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689
result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_cond,
result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689
result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689
result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689
result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_return_output);

-- t8_MUX_uxn_opcodes_h_l1416_c7_b689
t8_MUX_uxn_opcodes_h_l1416_c7_b689 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1416_c7_b689_cond,
t8_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue,
t8_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse,
t8_MUX_uxn_opcodes_h_l1416_c7_b689_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb
BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_left,
BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_right,
BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b
tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond,
tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue,
tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse,
tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b
result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond,
result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b
result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b
result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b
result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output);

-- t8_MUX_uxn_opcodes_h_l1419_c7_fa4b
t8_MUX_uxn_opcodes_h_l1419_c7_fa4b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond,
t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue,
t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse,
t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b
sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_ins,
sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_x,
sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_y,
sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3
BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3_left,
BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3_right,
BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1425_c7_7691
tmp8_MUX_uxn_opcodes_h_l1425_c7_7691 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_cond,
tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue,
tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse,
tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691
result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_cond,
result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691
result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691
result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691
result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b
BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b_left,
BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b_right,
BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75
tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_cond,
tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue,
tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse,
tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75
result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75
result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75
result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_cond,
result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1434_c11_6cab
BIN_OP_EQ_uxn_opcodes_h_l1434_c11_6cab : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1434_c11_6cab_left,
BIN_OP_EQ_uxn_opcodes_h_l1434_c11_6cab_right,
BIN_OP_EQ_uxn_opcodes_h_l1434_c11_6cab_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420
result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420
result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_return_output,
 tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output,
 t8_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_return_output,
 tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_return_output,
 t8_MUX_uxn_opcodes_h_l1416_c7_b689_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_return_output,
 tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output,
 t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output,
 sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3_return_output,
 tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b_return_output,
 tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1434_c11_6cab_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1413_c3_b6af : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1416_c7_b689_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1409_c2_b22e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1417_c3_0514 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1416_c7_b689_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1423_c22_fc1b_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1426_c3_6c95 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1431_c3_d126 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1434_c11_6cab_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1434_c11_6cab_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1434_c11_6cab_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1416_l1409_l1419_DUPLICATE_c7f8_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1409_l1428_l1425_l1419_l1416_DUPLICATE_3c98_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1409_l1434_l1425_l1419_l1416_DUPLICATE_8f90_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1425_l1416_l1409_DUPLICATE_d27d_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1434_l1428_l1425_l1419_l1416_DUPLICATE_d44f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1425_l1428_l1419_DUPLICATE_c483_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e78e_uxn_opcodes_h_l1439_l1405_DUPLICATE_9a75_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1434_c11_6cab_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1413_c3_b6af := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1413_c3_b6af;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1417_c3_0514 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1417_c3_0514;
     VAR_sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1426_c3_6c95 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1426_c3_6c95;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1431_c3_d126 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1431_c3_d126;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1434_c11_6cab_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse := tmp8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1428_c11_ba0b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1416_l1409_l1419_DUPLICATE_c7f8 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1416_l1409_l1419_DUPLICATE_c7f8_return_output := result.u16_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1434_l1428_l1425_l1419_l1416_DUPLICATE_d44f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1434_l1428_l1425_l1419_l1416_DUPLICATE_d44f_return_output := result.is_opc_done;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1423_c22_fc1b] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1423_c22_fc1b_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l1419_c11_a6bb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_left;
     BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_return_output := BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1425_l1416_l1409_DUPLICATE_d27d LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1425_l1416_l1409_DUPLICATE_d27d_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1425_l1428_l1419_DUPLICATE_c483 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1425_l1428_l1419_DUPLICATE_c483_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1434_c11_6cab] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1434_c11_6cab_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1434_c11_6cab_left;
     BIN_OP_EQ_uxn_opcodes_h_l1434_c11_6cab_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1434_c11_6cab_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1434_c11_6cab_return_output := BIN_OP_EQ_uxn_opcodes_h_l1434_c11_6cab_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1422_c30_c99b] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_ins;
     sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_x;
     sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_return_output := sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1416_c11_2f58] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_left;
     BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_return_output := BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1409_l1428_l1425_l1419_l1416_DUPLICATE_3c98 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1409_l1428_l1425_l1419_l1416_DUPLICATE_3c98_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1409_c6_4d0f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1409_l1434_l1425_l1419_l1416_DUPLICATE_8f90 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1409_l1434_l1425_l1419_l1416_DUPLICATE_8f90_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1425_c11_72a3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3_left;
     BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3_return_output := BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1409_c2_b22e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1409_c6_4d0f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1416_c7_b689_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1416_c11_2f58_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1419_c11_a6bb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1425_c11_72a3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1428_c11_ba0b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1434_c11_6cab_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1434_c11_6cab_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1423_c22_fc1b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1425_l1416_l1409_DUPLICATE_d27d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1425_l1416_l1409_DUPLICATE_d27d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1425_l1416_l1409_DUPLICATE_d27d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1416_l1409_l1419_DUPLICATE_c7f8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1416_l1409_l1419_DUPLICATE_c7f8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1416_l1409_l1419_DUPLICATE_c7f8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1434_l1428_l1425_l1419_l1416_DUPLICATE_d44f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1434_l1428_l1425_l1419_l1416_DUPLICATE_d44f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1434_l1428_l1425_l1419_l1416_DUPLICATE_d44f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1434_l1428_l1425_l1419_l1416_DUPLICATE_d44f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1434_l1428_l1425_l1419_l1416_DUPLICATE_d44f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1409_l1434_l1425_l1419_l1416_DUPLICATE_8f90_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1409_l1434_l1425_l1419_l1416_DUPLICATE_8f90_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1409_l1434_l1425_l1419_l1416_DUPLICATE_8f90_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1409_l1434_l1425_l1419_l1416_DUPLICATE_8f90_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1409_l1434_l1425_l1419_l1416_DUPLICATE_8f90_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1425_l1428_l1419_DUPLICATE_c483_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1425_l1428_l1419_DUPLICATE_c483_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1425_l1428_l1419_DUPLICATE_c483_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1409_l1428_l1425_l1419_l1416_DUPLICATE_3c98_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1409_l1428_l1425_l1419_l1416_DUPLICATE_3c98_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1409_l1428_l1425_l1419_l1416_DUPLICATE_3c98_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1409_l1428_l1425_l1419_l1416_DUPLICATE_3c98_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1409_l1428_l1425_l1419_l1416_DUPLICATE_3c98_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1422_c30_c99b_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1428_c7_ad75] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output;

     -- t8_MUX[uxn_opcodes_h_l1419_c7_fa4b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond <= VAR_t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond;
     t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue;
     t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output := t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1434_c7_9420] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1425_c7_7691] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1428_c7_ad75] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output := result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1419_c7_fa4b] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output := result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1428_c7_ad75] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_cond;
     tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output := tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1434_c7_9420] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1434_c7_9420_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1434_c7_9420_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1425_c7_7691_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1425_c7_7691] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_return_output;

     -- t8_MUX[uxn_opcodes_h_l1416_c7_b689] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1416_c7_b689_cond <= VAR_t8_MUX_uxn_opcodes_h_l1416_c7_b689_cond;
     t8_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue;
     t8_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1416_c7_b689_return_output := t8_MUX_uxn_opcodes_h_l1416_c7_b689_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1428_c7_ad75] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1419_c7_fa4b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1425_c7_7691] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_return_output := result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1425_c7_7691] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_cond;
     tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_return_output := tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1416_c7_b689] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_return_output := result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1428_c7_ad75] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1428_c7_ad75_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1425_c7_7691_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1416_c7_b689_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1425_c7_7691_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1416_c7_b689_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1425_c7_7691_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1425_c7_7691] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1419_c7_fa4b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output;

     -- t8_MUX[uxn_opcodes_h_l1409_c2_b22e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1409_c2_b22e_cond <= VAR_t8_MUX_uxn_opcodes_h_l1409_c2_b22e_cond;
     t8_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue;
     t8_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output := t8_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1416_c7_b689] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1419_c7_fa4b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1419_c7_fa4b] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond;
     tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output := tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1425_c7_7691] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1409_c2_b22e] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output := result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1425_c7_7691_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1425_c7_7691_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1416_c7_b689_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1419_c7_fa4b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1409_c2_b22e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1416_c7_b689] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_return_output := result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1416_c7_b689] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1416_c7_b689] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_cond;
     tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_return_output := tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1419_c7_fa4b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1419_c7_fa4b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1416_c7_b689_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1416_c7_b689_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1416_c7_b689_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1416_c7_b689] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1416_c7_b689] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1409_c2_b22e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1409_c2_b22e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output := result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1409_c2_b22e] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_cond;
     tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output := tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1416_c7_b689_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1416_c7_b689_return_output;
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1409_c2_b22e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1409_c2_b22e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_e78e_uxn_opcodes_h_l1439_l1405_DUPLICATE_9a75 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e78e_uxn_opcodes_h_l1439_l1405_DUPLICATE_9a75_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_e78e(
     result,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1409_c2_b22e_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e78e_uxn_opcodes_h_l1439_l1405_DUPLICATE_9a75_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e78e_uxn_opcodes_h_l1439_l1405_DUPLICATE_9a75_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
