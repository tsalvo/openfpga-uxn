-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 37
entity nip_0CLK_d7ba9283 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end nip_0CLK_d7ba9283;
architecture arch of nip_0CLK_d7ba9283 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2333_c6_c5bd]
signal BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2333_c2_ed12]
signal t8_MUX_uxn_opcodes_h_l2333_c2_ed12_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2333_c2_ed12]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2333_c2_ed12]
signal result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2333_c2_ed12]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2333_c2_ed12]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2333_c2_ed12]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2333_c2_ed12]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2338_c11_185b]
signal BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2338_c7_4f29]
signal t8_MUX_uxn_opcodes_h_l2338_c7_4f29_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2338_c7_4f29]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2338_c7_4f29]
signal result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2338_c7_4f29]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2338_c7_4f29]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2338_c7_4f29]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2338_c7_4f29]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2341_c11_dc30]
signal BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2341_c7_c12b]
signal t8_MUX_uxn_opcodes_h_l2341_c7_c12b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2341_c7_c12b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2341_c7_c12b]
signal result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2341_c7_c12b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2341_c7_c12b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2341_c7_c12b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2341_c7_c12b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l2344_c32_988b]
signal BIN_OP_AND_uxn_opcodes_h_l2344_c32_988b_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2344_c32_988b_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2344_c32_988b_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l2344_c32_45e7]
signal BIN_OP_GT_uxn_opcodes_h_l2344_c32_45e7_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l2344_c32_45e7_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l2344_c32_45e7_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l2344_c32_3a81]
signal MUX_uxn_opcodes_h_l2344_c32_3a81_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l2344_c32_3a81_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l2344_c32_3a81_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l2344_c32_3a81_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2346_c11_35db]
signal BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2346_c7_3dab]
signal result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2346_c7_3dab]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2346_c7_3dab]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2346_c7_3dab]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2346_c7_3dab]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2352_c11_1208]
signal BIN_OP_EQ_uxn_opcodes_h_l2352_c11_1208_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2352_c11_1208_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2352_c11_1208_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2352_c7_9bac]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2352_c7_9bac]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_value := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_sp_shift := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.is_opc_done := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd
BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_left,
BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_right,
BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_return_output);

-- t8_MUX_uxn_opcodes_h_l2333_c2_ed12
t8_MUX_uxn_opcodes_h_l2333_c2_ed12 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2333_c2_ed12_cond,
t8_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue,
t8_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse,
t8_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12
result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12
result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_cond,
result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12
result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12
result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12
result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b
BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_left,
BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_right,
BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_return_output);

-- t8_MUX_uxn_opcodes_h_l2338_c7_4f29
t8_MUX_uxn_opcodes_h_l2338_c7_4f29 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2338_c7_4f29_cond,
t8_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue,
t8_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse,
t8_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29
result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29
result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_cond,
result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29
result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29
result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29
result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30
BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_left,
BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_right,
BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_return_output);

-- t8_MUX_uxn_opcodes_h_l2341_c7_c12b
t8_MUX_uxn_opcodes_h_l2341_c7_c12b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2341_c7_c12b_cond,
t8_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue,
t8_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse,
t8_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b
result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b
result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_cond,
result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b
result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b
result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b
result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l2344_c32_988b
BIN_OP_AND_uxn_opcodes_h_l2344_c32_988b : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l2344_c32_988b_left,
BIN_OP_AND_uxn_opcodes_h_l2344_c32_988b_right,
BIN_OP_AND_uxn_opcodes_h_l2344_c32_988b_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l2344_c32_45e7
BIN_OP_GT_uxn_opcodes_h_l2344_c32_45e7 : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l2344_c32_45e7_left,
BIN_OP_GT_uxn_opcodes_h_l2344_c32_45e7_right,
BIN_OP_GT_uxn_opcodes_h_l2344_c32_45e7_return_output);

-- MUX_uxn_opcodes_h_l2344_c32_3a81
MUX_uxn_opcodes_h_l2344_c32_3a81 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l2344_c32_3a81_cond,
MUX_uxn_opcodes_h_l2344_c32_3a81_iftrue,
MUX_uxn_opcodes_h_l2344_c32_3a81_iffalse,
MUX_uxn_opcodes_h_l2344_c32_3a81_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db
BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db_left,
BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db_right,
BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab
result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_cond,
result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab
result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab
result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab
result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2352_c11_1208
BIN_OP_EQ_uxn_opcodes_h_l2352_c11_1208 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2352_c11_1208_left,
BIN_OP_EQ_uxn_opcodes_h_l2352_c11_1208_right,
BIN_OP_EQ_uxn_opcodes_h_l2352_c11_1208_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac
result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac
result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_return_output,
 t8_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_return_output,
 t8_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_return_output,
 t8_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output,
 BIN_OP_AND_uxn_opcodes_h_l2344_c32_988b_return_output,
 BIN_OP_GT_uxn_opcodes_h_l2344_c32_45e7_return_output,
 MUX_uxn_opcodes_h_l2344_c32_3a81_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2352_c11_1208_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2333_c2_ed12_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2335_c3_dba7 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2338_c7_4f29_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2339_c3_314a : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2341_c7_c12b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2344_c32_3a81_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2344_c32_3a81_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2344_c32_3a81_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2344_c32_988b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2344_c32_988b_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2344_c32_988b_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2344_c32_45e7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2344_c32_45e7_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2344_c32_45e7_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2344_c32_3a81_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2349_c3_b57c : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_1208_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_1208_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_1208_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2341_l2333_l2338_DUPLICATE_2c46_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2341_l2333_l2346_l2338_DUPLICATE_968b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2333_l2346_l2338_DUPLICATE_5d6f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2352_l2341_l2333_l2338_DUPLICATE_e5fb_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2352_l2341_l2346_l2338_DUPLICATE_0348_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2341_l2346_DUPLICATE_f224_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l2357_l2329_DUPLICATE_a35e_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db_right := to_unsigned(3, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l2344_c32_3a81_iftrue := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l2344_c32_3a81_iffalse := resize(to_signed(-1, 2), 8);
     VAR_BIN_OP_AND_uxn_opcodes_h_l2344_c32_988b_right := to_unsigned(128, 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2349_c3_b57c := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2349_c3_b57c;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2339_c3_314a := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2339_c3_314a;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2335_c3_dba7 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2335_c3_dba7;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_1208_right := to_unsigned(4, 3);
     VAR_BIN_OP_GT_uxn_opcodes_h_l2344_c32_45e7_right := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_right := to_unsigned(2, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_BIN_OP_AND_uxn_opcodes_h_l2344_c32_988b_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_1208_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue := VAR_previous_stack_read;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2338_c11_185b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_left;
     BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_return_output := BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_return_output;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2341_l2333_l2338_DUPLICATE_2c46 LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2341_l2333_l2338_DUPLICATE_2c46_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2352_l2341_l2346_l2338_DUPLICATE_0348 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2352_l2341_l2346_l2338_DUPLICATE_0348_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2333_c6_c5bd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_left;
     BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_return_output := BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2352_l2341_l2333_l2338_DUPLICATE_e5fb LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2352_l2341_l2333_l2338_DUPLICATE_e5fb_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2341_l2333_l2346_l2338_DUPLICATE_968b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2341_l2333_l2346_l2338_DUPLICATE_968b_return_output := result.stack_value;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2341_l2346_DUPLICATE_f224 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2341_l2346_DUPLICATE_f224_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2352_c11_1208] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2352_c11_1208_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_1208_left;
     BIN_OP_EQ_uxn_opcodes_h_l2352_c11_1208_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_1208_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_1208_return_output := BIN_OP_EQ_uxn_opcodes_h_l2352_c11_1208_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2333_l2346_l2338_DUPLICATE_5d6f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2333_l2346_l2338_DUPLICATE_5d6f_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2346_c11_35db] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db_left;
     BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db_return_output := BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2341_c11_dc30] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_left;
     BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_return_output := BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l2344_c32_988b] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l2344_c32_988b_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l2344_c32_988b_left;
     BIN_OP_AND_uxn_opcodes_h_l2344_c32_988b_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l2344_c32_988b_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l2344_c32_988b_return_output := BIN_OP_AND_uxn_opcodes_h_l2344_c32_988b_return_output;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l2344_c32_45e7_left := VAR_BIN_OP_AND_uxn_opcodes_h_l2344_c32_988b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2333_c2_ed12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2333_c6_c5bd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2338_c7_4f29_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2338_c11_185b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2341_c7_c12b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2341_c11_dc30_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_35db_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_1208_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2352_c11_1208_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2341_l2333_l2338_DUPLICATE_2c46_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2341_l2333_l2338_DUPLICATE_2c46_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2341_l2333_l2338_DUPLICATE_2c46_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2352_l2341_l2346_l2338_DUPLICATE_0348_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2352_l2341_l2346_l2338_DUPLICATE_0348_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2352_l2341_l2346_l2338_DUPLICATE_0348_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2352_l2341_l2346_l2338_DUPLICATE_0348_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2333_l2346_l2338_DUPLICATE_5d6f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2333_l2346_l2338_DUPLICATE_5d6f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2333_l2346_l2338_DUPLICATE_5d6f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2352_l2341_l2333_l2338_DUPLICATE_e5fb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2352_l2341_l2333_l2338_DUPLICATE_e5fb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2352_l2341_l2333_l2338_DUPLICATE_e5fb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2352_l2341_l2333_l2338_DUPLICATE_e5fb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2341_l2346_DUPLICATE_f224_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2341_l2346_DUPLICATE_f224_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2341_l2333_l2346_l2338_DUPLICATE_968b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2341_l2333_l2346_l2338_DUPLICATE_968b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2341_l2333_l2346_l2338_DUPLICATE_968b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2341_l2333_l2346_l2338_DUPLICATE_968b_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2346_c7_3dab] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2346_c7_3dab] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l2344_c32_45e7] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l2344_c32_45e7_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l2344_c32_45e7_left;
     BIN_OP_GT_uxn_opcodes_h_l2344_c32_45e7_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l2344_c32_45e7_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l2344_c32_45e7_return_output := BIN_OP_GT_uxn_opcodes_h_l2344_c32_45e7_return_output;

     -- t8_MUX[uxn_opcodes_h_l2341_c7_c12b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2341_c7_c12b_cond <= VAR_t8_MUX_uxn_opcodes_h_l2341_c7_c12b_cond;
     t8_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue;
     t8_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output := t8_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2352_c7_9bac] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2352_c7_9bac] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2346_c7_3dab] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output := result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l2344_c32_3a81_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l2344_c32_45e7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2352_c7_9bac_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2352_c7_9bac_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2341_c7_c12b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output;

     -- MUX[uxn_opcodes_h_l2344_c32_3a81] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l2344_c32_3a81_cond <= VAR_MUX_uxn_opcodes_h_l2344_c32_3a81_cond;
     MUX_uxn_opcodes_h_l2344_c32_3a81_iftrue <= VAR_MUX_uxn_opcodes_h_l2344_c32_3a81_iftrue;
     MUX_uxn_opcodes_h_l2344_c32_3a81_iffalse <= VAR_MUX_uxn_opcodes_h_l2344_c32_3a81_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l2344_c32_3a81_return_output := MUX_uxn_opcodes_h_l2344_c32_3a81_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2346_c7_3dab] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output;

     -- t8_MUX[uxn_opcodes_h_l2338_c7_4f29] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2338_c7_4f29_cond <= VAR_t8_MUX_uxn_opcodes_h_l2338_c7_4f29_cond;
     t8_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue;
     t8_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output := t8_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2341_c7_c12b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2341_c7_c12b] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output := result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2346_c7_3dab] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue := VAR_MUX_uxn_opcodes_h_l2344_c32_3a81_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_3dab_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output;
     -- t8_MUX[uxn_opcodes_h_l2333_c2_ed12] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2333_c2_ed12_cond <= VAR_t8_MUX_uxn_opcodes_h_l2333_c2_ed12_cond;
     t8_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue;
     t8_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output := t8_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2341_c7_c12b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2338_c7_4f29] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output := result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2338_c7_4f29] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2341_c7_c12b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2338_c7_4f29] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2341_c7_c12b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2341_c7_c12b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2338_c7_4f29] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2338_c7_4f29] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2338_c7_4f29] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2333_c2_ed12] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2333_c2_ed12] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output := result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2333_c2_ed12] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2338_c7_4f29_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2333_c2_ed12] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2333_c2_ed12] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2333_c2_ed12] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l2357_l2329_DUPLICATE_a35e LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l2357_l2329_DUPLICATE_a35e_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2333_c2_ed12_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l2357_l2329_DUPLICATE_a35e_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l2357_l2329_DUPLICATE_a35e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
