-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity lth2_0CLK_85d5529e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(15 downto 0);
 return_output : out opcode_result_t);
end lth2_0CLK_85d5529e;
architecture arch of lth2_0CLK_85d5529e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1757_c6_a1e0]
signal BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1757_c2_1363]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1757_c2_1363]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1757_c2_1363]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1757_c2_1363]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1757_c2_1363]
signal result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1757_c2_1363]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1757_c2_1363]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l1757_c2_1363]
signal n16_MUX_uxn_opcodes_h_l1757_c2_1363_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1757_c2_1363_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l1757_c2_1363]
signal t16_MUX_uxn_opcodes_h_l1757_c2_1363_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1757_c2_1363_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1765_c11_0544]
signal BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1765_c7_3dc0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1765_c7_3dc0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1765_c7_3dc0]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1765_c7_3dc0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1765_c7_3dc0]
signal result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1765_c7_3dc0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1765_c7_3dc0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l1765_c7_3dc0]
signal n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l1765_c7_3dc0]
signal t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1768_c11_c459]
signal BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1768_c7_1cd0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1768_c7_1cd0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1768_c7_1cd0]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1768_c7_1cd0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1768_c7_1cd0]
signal result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1768_c7_1cd0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1768_c7_1cd0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l1768_c7_1cd0]
signal n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l1768_c7_1cd0]
signal t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1772_c30_abab]
signal sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1774_c11_f373]
signal BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1774_c7_a915]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1774_c7_a915]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1774_c7_a915]
signal result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1774_c7_a915]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1774_c7_a915]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_return_output : unsigned(3 downto 0);

-- n16_MUX[uxn_opcodes_h_l1774_c7_a915]
signal n16_MUX_uxn_opcodes_h_l1774_c7_a915_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1774_c7_a915_return_output : unsigned(15 downto 0);

-- BIN_OP_LT[uxn_opcodes_h_l1779_c21_0a88]
signal BIN_OP_LT_uxn_opcodes_h_l1779_c21_0a88_left : unsigned(15 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l1779_c21_0a88_right : unsigned(15 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l1779_c21_0a88_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1779_c21_80ab]
signal MUX_uxn_opcodes_h_l1779_c21_80ab_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1779_c21_80ab_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1779_c21_80ab_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1779_c21_80ab_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1781_c11_178f]
signal BIN_OP_EQ_uxn_opcodes_h_l1781_c11_178f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1781_c11_178f_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1781_c11_178f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1781_c7_ba60]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1781_c7_ba60]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_stack_operation_16bit := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_stack_write := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0
BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_left,
BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_right,
BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363
result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363
result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363
result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_cond,
result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363
result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363
result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_return_output);

-- n16_MUX_uxn_opcodes_h_l1757_c2_1363
n16_MUX_uxn_opcodes_h_l1757_c2_1363 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1757_c2_1363_cond,
n16_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue,
n16_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse,
n16_MUX_uxn_opcodes_h_l1757_c2_1363_return_output);

-- t16_MUX_uxn_opcodes_h_l1757_c2_1363
t16_MUX_uxn_opcodes_h_l1757_c2_1363 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1757_c2_1363_cond,
t16_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue,
t16_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse,
t16_MUX_uxn_opcodes_h_l1757_c2_1363_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544
BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_left,
BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_right,
BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0
result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0
result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0
result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond,
result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0
result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0
result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output);

-- n16_MUX_uxn_opcodes_h_l1765_c7_3dc0
n16_MUX_uxn_opcodes_h_l1765_c7_3dc0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond,
n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue,
n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse,
n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output);

-- t16_MUX_uxn_opcodes_h_l1765_c7_3dc0
t16_MUX_uxn_opcodes_h_l1765_c7_3dc0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond,
t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue,
t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse,
t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459
BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_left,
BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_right,
BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0
result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0
result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0
result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond,
result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0
result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0
result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output);

-- n16_MUX_uxn_opcodes_h_l1768_c7_1cd0
n16_MUX_uxn_opcodes_h_l1768_c7_1cd0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond,
n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue,
n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse,
n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output);

-- t16_MUX_uxn_opcodes_h_l1768_c7_1cd0
t16_MUX_uxn_opcodes_h_l1768_c7_1cd0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond,
t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue,
t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse,
t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1772_c30_abab
sp_relative_shift_uxn_opcodes_h_l1772_c30_abab : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_ins,
sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_x,
sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_y,
sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373
BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373_left,
BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373_right,
BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915
result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915
result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915
result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_cond,
result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915
result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_return_output);

-- n16_MUX_uxn_opcodes_h_l1774_c7_a915
n16_MUX_uxn_opcodes_h_l1774_c7_a915 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1774_c7_a915_cond,
n16_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue,
n16_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse,
n16_MUX_uxn_opcodes_h_l1774_c7_a915_return_output);

-- BIN_OP_LT_uxn_opcodes_h_l1779_c21_0a88
BIN_OP_LT_uxn_opcodes_h_l1779_c21_0a88 : entity work.BIN_OP_LT_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_LT_uxn_opcodes_h_l1779_c21_0a88_left,
BIN_OP_LT_uxn_opcodes_h_l1779_c21_0a88_right,
BIN_OP_LT_uxn_opcodes_h_l1779_c21_0a88_return_output);

-- MUX_uxn_opcodes_h_l1779_c21_80ab
MUX_uxn_opcodes_h_l1779_c21_80ab : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1779_c21_80ab_cond,
MUX_uxn_opcodes_h_l1779_c21_80ab_iftrue,
MUX_uxn_opcodes_h_l1779_c21_80ab_iffalse,
MUX_uxn_opcodes_h_l1779_c21_80ab_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1781_c11_178f
BIN_OP_EQ_uxn_opcodes_h_l1781_c11_178f : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1781_c11_178f_left,
BIN_OP_EQ_uxn_opcodes_h_l1781_c11_178f_right,
BIN_OP_EQ_uxn_opcodes_h_l1781_c11_178f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60
result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60
result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_return_output,
 n16_MUX_uxn_opcodes_h_l1757_c2_1363_return_output,
 t16_MUX_uxn_opcodes_h_l1757_c2_1363_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output,
 n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output,
 t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output,
 n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output,
 t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output,
 sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_return_output,
 n16_MUX_uxn_opcodes_h_l1774_c7_a915_return_output,
 BIN_OP_LT_uxn_opcodes_h_l1779_c21_0a88_return_output,
 MUX_uxn_opcodes_h_l1779_c21_80ab_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1781_c11_178f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1762_c3_288c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1757_c2_1363_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1757_c2_1363_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1757_c2_1363_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1757_c2_1363_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1766_c3_a293 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1774_c7_a915_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1778_c3_9de4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1774_c7_a915_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1779_c21_80ab_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1779_c21_0a88_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1779_c21_0a88_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1779_c21_0a88_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1779_c21_80ab_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1779_c21_80ab_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1779_c21_80ab_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1781_c11_178f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1781_c11_178f_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1781_c11_178f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1774_l1765_l1757_DUPLICATE_ae0e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1774_l1765_l1768_l1757_DUPLICATE_5f4c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1765_l1768_l1757_DUPLICATE_0dc8_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1765_l1781_l1768_l1757_DUPLICATE_7335_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1765_l1768_DUPLICATE_e3db_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1774_l1765_l1781_l1768_DUPLICATE_2db5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1774_l1768_DUPLICATE_d598_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a_uxn_opcodes_h_l1786_l1753_DUPLICATE_24b7_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n16 := n16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_MUX_uxn_opcodes_h_l1779_c21_80ab_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1778_c3_9de4 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1778_c3_9de4;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1766_c3_a293 := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1766_c3_a293;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_y := resize(to_signed(-3, 3), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1781_c11_178f_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1762_c3_288c := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1762_c3_288c;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_right := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1779_c21_80ab_iftrue := resize(to_unsigned(1, 1), 8);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_ins := VAR_ins;
     VAR_n16_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse := n16;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1781_c11_178f_left := VAR_phase;
     VAR_BIN_OP_LT_uxn_opcodes_h_l1779_c21_0a88_left := VAR_previous_stack_read;
     VAR_n16_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue := VAR_previous_stack_read;
     VAR_t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_LT_uxn_opcodes_h_l1779_c21_0a88_right := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse := t16;
     -- BIN_OP_EQ[uxn_opcodes_h_l1781_c11_178f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1781_c11_178f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1781_c11_178f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1781_c11_178f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1781_c11_178f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1781_c11_178f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1781_c11_178f_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1774_l1765_l1768_l1757_DUPLICATE_5f4c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1774_l1765_l1768_l1757_DUPLICATE_5f4c_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1774_l1765_l1781_l1768_DUPLICATE_2db5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1774_l1765_l1781_l1768_DUPLICATE_2db5_return_output := result.is_opc_done;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1765_l1768_l1757_DUPLICATE_0dc8 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1765_l1768_l1757_DUPLICATE_0dc8_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1765_c11_0544] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_left;
     BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_return_output := BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1765_l1768_DUPLICATE_e3db LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1765_l1768_DUPLICATE_e3db_return_output := result.is_stack_operation_16bit;

     -- BIN_OP_LT[uxn_opcodes_h_l1779_c21_0a88] LATENCY=0
     -- Inputs
     BIN_OP_LT_uxn_opcodes_h_l1779_c21_0a88_left <= VAR_BIN_OP_LT_uxn_opcodes_h_l1779_c21_0a88_left;
     BIN_OP_LT_uxn_opcodes_h_l1779_c21_0a88_right <= VAR_BIN_OP_LT_uxn_opcodes_h_l1779_c21_0a88_right;
     -- Outputs
     VAR_BIN_OP_LT_uxn_opcodes_h_l1779_c21_0a88_return_output := BIN_OP_LT_uxn_opcodes_h_l1779_c21_0a88_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1774_l1768_DUPLICATE_d598 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1774_l1768_DUPLICATE_d598_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1768_c11_c459] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_left;
     BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_return_output := BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1757_c6_a1e0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_left;
     BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_return_output := BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1774_c11_f373] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373_left;
     BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373_return_output := BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1772_c30_abab] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_ins;
     sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_x;
     sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_return_output := sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1765_l1781_l1768_l1757_DUPLICATE_7335 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1765_l1781_l1768_l1757_DUPLICATE_7335_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1774_l1765_l1757_DUPLICATE_ae0e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1774_l1765_l1757_DUPLICATE_ae0e_return_output := result.is_sp_shift;

     -- Submodule level 1
     VAR_n16_MUX_uxn_opcodes_h_l1757_c2_1363_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1757_c2_1363_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1757_c6_a1e0_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1765_c11_0544_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1768_c11_c459_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1774_c7_a915_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1774_c11_f373_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1781_c11_178f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1781_c11_178f_return_output;
     VAR_MUX_uxn_opcodes_h_l1779_c21_80ab_cond := VAR_BIN_OP_LT_uxn_opcodes_h_l1779_c21_0a88_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1765_l1768_l1757_DUPLICATE_0dc8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1765_l1768_l1757_DUPLICATE_0dc8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1765_l1768_l1757_DUPLICATE_0dc8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1774_l1765_l1781_l1768_DUPLICATE_2db5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1774_l1765_l1781_l1768_DUPLICATE_2db5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1774_l1765_l1781_l1768_DUPLICATE_2db5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1774_l1765_l1781_l1768_DUPLICATE_2db5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1774_l1765_l1757_DUPLICATE_ae0e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1774_l1765_l1757_DUPLICATE_ae0e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1774_l1765_l1757_DUPLICATE_ae0e_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1765_l1768_DUPLICATE_e3db_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1765_l1768_DUPLICATE_e3db_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1765_l1781_l1768_l1757_DUPLICATE_7335_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1765_l1781_l1768_l1757_DUPLICATE_7335_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1765_l1781_l1768_l1757_DUPLICATE_7335_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1765_l1781_l1768_l1757_DUPLICATE_7335_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1774_l1768_DUPLICATE_d598_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1774_l1768_DUPLICATE_d598_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1774_l1765_l1768_l1757_DUPLICATE_5f4c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1774_l1765_l1768_l1757_DUPLICATE_5f4c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1774_l1765_l1768_l1757_DUPLICATE_5f4c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1774_l1765_l1768_l1757_DUPLICATE_5f4c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1772_c30_abab_return_output;
     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1768_c7_1cd0] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1774_c7_a915] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_return_output;

     -- n16_MUX[uxn_opcodes_h_l1774_c7_a915] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1774_c7_a915_cond <= VAR_n16_MUX_uxn_opcodes_h_l1774_c7_a915_cond;
     n16_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue;
     n16_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1774_c7_a915_return_output := n16_MUX_uxn_opcodes_h_l1774_c7_a915_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1781_c7_ba60] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1774_c7_a915] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_return_output;

     -- MUX[uxn_opcodes_h_l1779_c21_80ab] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1779_c21_80ab_cond <= VAR_MUX_uxn_opcodes_h_l1779_c21_80ab_cond;
     MUX_uxn_opcodes_h_l1779_c21_80ab_iftrue <= VAR_MUX_uxn_opcodes_h_l1779_c21_80ab_iftrue;
     MUX_uxn_opcodes_h_l1779_c21_80ab_iffalse <= VAR_MUX_uxn_opcodes_h_l1779_c21_80ab_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1779_c21_80ab_return_output := MUX_uxn_opcodes_h_l1779_c21_80ab_return_output;

     -- t16_MUX[uxn_opcodes_h_l1768_c7_1cd0] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond <= VAR_t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond;
     t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue;
     t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output := t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1768_c7_1cd0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1781_c7_ba60] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue := VAR_MUX_uxn_opcodes_h_l1779_c21_80ab_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1774_c7_a915_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1781_c7_ba60_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1774_c7_a915_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1781_c7_ba60_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1774_c7_a915_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output;
     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1765_c7_3dc0] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1765_c7_3dc0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1768_c7_1cd0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1768_c7_1cd0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1774_c7_a915] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_return_output;

     -- n16_MUX[uxn_opcodes_h_l1768_c7_1cd0] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond <= VAR_n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond;
     n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue;
     n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output := n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1774_c7_a915] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_return_output;

     -- t16_MUX[uxn_opcodes_h_l1765_c7_3dc0] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond <= VAR_t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond;
     t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue;
     t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output := t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1774_c7_a915] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_return_output := result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_return_output;

     -- Submodule level 3
     VAR_n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1774_c7_a915_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1774_c7_a915_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1774_c7_a915_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1765_c7_3dc0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output;

     -- t16_MUX[uxn_opcodes_h_l1757_c2_1363] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1757_c2_1363_cond <= VAR_t16_MUX_uxn_opcodes_h_l1757_c2_1363_cond;
     t16_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue;
     t16_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1757_c2_1363_return_output := t16_MUX_uxn_opcodes_h_l1757_c2_1363_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1768_c7_1cd0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output := result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1768_c7_1cd0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1757_c2_1363] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_return_output;

     -- n16_MUX[uxn_opcodes_h_l1765_c7_3dc0] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond <= VAR_n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond;
     n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue;
     n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output := n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1765_c7_3dc0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1757_c2_1363] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1768_c7_1cd0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output;

     -- Submodule level 4
     VAR_n16_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1768_c7_1cd0_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l1757_c2_1363_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1765_c7_3dc0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1757_c2_1363] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1757_c2_1363] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1765_c7_3dc0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output;

     -- n16_MUX[uxn_opcodes_h_l1757_c2_1363] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1757_c2_1363_cond <= VAR_n16_MUX_uxn_opcodes_h_l1757_c2_1363_cond;
     n16_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue;
     n16_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1757_c2_1363_return_output := n16_MUX_uxn_opcodes_h_l1757_c2_1363_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1765_c7_3dc0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output := result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output;

     -- Submodule level 5
     REG_VAR_n16 := VAR_n16_MUX_uxn_opcodes_h_l1757_c2_1363_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1765_c7_3dc0_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1757_c2_1363] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1757_c2_1363] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1757_c2_1363] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_return_output := result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a_uxn_opcodes_h_l1786_l1753_DUPLICATE_24b7 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a_uxn_opcodes_h_l1786_l1753_DUPLICATE_24b7_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1757_c2_1363_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1757_c2_1363_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1757_c2_1363_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1757_c2_1363_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1757_c2_1363_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1757_c2_1363_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1757_c2_1363_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a_uxn_opcodes_h_l1786_l1753_DUPLICATE_24b7_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a_uxn_opcodes_h_l1786_l1753_DUPLICATE_24b7_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n16 <= REG_VAR_n16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n16 <= REG_COMB_n16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
