-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity neq_0CLK_7883ef49 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end neq_0CLK_7883ef49;
architecture arch of neq_0CLK_7883ef49 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1218_c6_7b8d]
signal BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1218_c2_4baf]
signal n8_MUX_uxn_opcodes_h_l1218_c2_4baf_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1218_c2_4baf]
signal result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1218_c2_4baf]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1218_c2_4baf]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1218_c2_4baf]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1218_c2_4baf]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1218_c2_4baf]
signal t8_MUX_uxn_opcodes_h_l1218_c2_4baf_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1225_c11_2770]
signal BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1225_c7_477a]
signal n8_MUX_uxn_opcodes_h_l1225_c7_477a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1225_c7_477a_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1225_c7_477a]
signal result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1225_c7_477a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1225_c7_477a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1225_c7_477a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1225_c7_477a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1225_c7_477a]
signal t8_MUX_uxn_opcodes_h_l1225_c7_477a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1225_c7_477a_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1228_c11_fcc6]
signal BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1228_c7_ac0c]
signal n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1228_c7_ac0c]
signal result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1228_c7_ac0c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1228_c7_ac0c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1228_c7_ac0c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1228_c7_ac0c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1228_c7_ac0c]
signal t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1231_c11_8493]
signal BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1231_c7_5bf9]
signal n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1231_c7_5bf9]
signal result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1231_c7_5bf9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1231_c7_5bf9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1231_c7_5bf9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1231_c7_5bf9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output : signed(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1234_c30_ed5a]
signal sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1237_c21_c1f1]
signal BIN_OP_EQ_uxn_opcodes_h_l1237_c21_c1f1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1237_c21_c1f1_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1237_c21_c1f1_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1237_c21_e026]
signal MUX_uxn_opcodes_h_l1237_c21_e026_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1237_c21_e026_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1237_c21_e026_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1237_c21_e026_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1239_c11_624d]
signal BIN_OP_EQ_uxn_opcodes_h_l1239_c11_624d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1239_c11_624d_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1239_c11_624d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1239_c7_ddaa]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1239_c7_ddaa]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1239_c7_ddaa]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_return_output : signed(3 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_eae7( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.stack_address_sp_offset := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d
BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_left,
BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_right,
BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_return_output);

-- n8_MUX_uxn_opcodes_h_l1218_c2_4baf
n8_MUX_uxn_opcodes_h_l1218_c2_4baf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1218_c2_4baf_cond,
n8_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue,
n8_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse,
n8_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf
result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_cond,
result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf
result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf
result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf
result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output);

-- t8_MUX_uxn_opcodes_h_l1218_c2_4baf
t8_MUX_uxn_opcodes_h_l1218_c2_4baf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1218_c2_4baf_cond,
t8_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue,
t8_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse,
t8_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770
BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_left,
BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_right,
BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_return_output);

-- n8_MUX_uxn_opcodes_h_l1225_c7_477a
n8_MUX_uxn_opcodes_h_l1225_c7_477a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1225_c7_477a_cond,
n8_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue,
n8_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse,
n8_MUX_uxn_opcodes_h_l1225_c7_477a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a
result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_cond,
result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a
result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a
result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a
result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_return_output);

-- t8_MUX_uxn_opcodes_h_l1225_c7_477a
t8_MUX_uxn_opcodes_h_l1225_c7_477a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1225_c7_477a_cond,
t8_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue,
t8_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse,
t8_MUX_uxn_opcodes_h_l1225_c7_477a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6
BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_left,
BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_right,
BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_return_output);

-- n8_MUX_uxn_opcodes_h_l1228_c7_ac0c
n8_MUX_uxn_opcodes_h_l1228_c7_ac0c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond,
n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue,
n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse,
n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c
result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c
result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c
result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c
result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output);

-- t8_MUX_uxn_opcodes_h_l1228_c7_ac0c
t8_MUX_uxn_opcodes_h_l1228_c7_ac0c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond,
t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue,
t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse,
t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493
BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493_left,
BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493_right,
BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493_return_output);

-- n8_MUX_uxn_opcodes_h_l1231_c7_5bf9
n8_MUX_uxn_opcodes_h_l1231_c7_5bf9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond,
n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue,
n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse,
n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9
result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond,
result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9
result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9
result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9
result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a
sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_ins,
sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_x,
sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_y,
sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1237_c21_c1f1
BIN_OP_EQ_uxn_opcodes_h_l1237_c21_c1f1 : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1237_c21_c1f1_left,
BIN_OP_EQ_uxn_opcodes_h_l1237_c21_c1f1_right,
BIN_OP_EQ_uxn_opcodes_h_l1237_c21_c1f1_return_output);

-- MUX_uxn_opcodes_h_l1237_c21_e026
MUX_uxn_opcodes_h_l1237_c21_e026 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1237_c21_e026_cond,
MUX_uxn_opcodes_h_l1237_c21_e026_iftrue,
MUX_uxn_opcodes_h_l1237_c21_e026_iffalse,
MUX_uxn_opcodes_h_l1237_c21_e026_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1239_c11_624d
BIN_OP_EQ_uxn_opcodes_h_l1239_c11_624d : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1239_c11_624d_left,
BIN_OP_EQ_uxn_opcodes_h_l1239_c11_624d_right,
BIN_OP_EQ_uxn_opcodes_h_l1239_c11_624d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa
result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa
result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa
result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_return_output,
 n8_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output,
 t8_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_return_output,
 n8_MUX_uxn_opcodes_h_l1225_c7_477a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_return_output,
 t8_MUX_uxn_opcodes_h_l1225_c7_477a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_return_output,
 n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output,
 t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493_return_output,
 n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output,
 sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1237_c21_c1f1_return_output,
 MUX_uxn_opcodes_h_l1237_c21_e026_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1239_c11_624d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1225_c7_477a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1218_c2_4baf_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1222_c3_eeed : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1225_c7_477a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1218_c2_4baf_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1225_c7_477a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1226_c3_a4cf : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1225_c7_477a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1236_c3_04ad : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1237_c21_e026_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c21_c1f1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c21_c1f1_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c21_c1f1_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1237_c21_e026_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1237_c21_e026_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1237_c21_e026_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_624d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_624d_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_624d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1240_c3_ebb4 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1218_l1225_l1228_l1231_DUPLICATE_2373_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1218_l1225_l1228_l1239_DUPLICATE_bbcd_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1218_l1225_l1228_l1239_DUPLICATE_1934_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1239_l1225_l1228_l1231_DUPLICATE_0679_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1228_l1231_DUPLICATE_b093_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1214_l1245_DUPLICATE_ab89_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493_right := to_unsigned(3, 2);
     VAR_MUX_uxn_opcodes_h_l1237_c21_e026_iffalse := resize(to_unsigned(1, 1), 8);
     VAR_MUX_uxn_opcodes_h_l1237_c21_e026_iftrue := resize(to_unsigned(0, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1222_c3_eeed := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1222_c3_eeed;
     VAR_sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1236_c3_04ad := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1236_c3_04ad;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_624d_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1226_c3_a4cf := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1226_c3_a4cf;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_right := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1240_c3_ebb4 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1240_c3_ebb4;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_624d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c21_c1f1_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c21_c1f1_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1225_c11_2770] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_left;
     BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_return_output := BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1239_l1225_l1228_l1231_DUPLICATE_0679 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1239_l1225_l1228_l1231_DUPLICATE_0679_return_output := result.is_opc_done;

     -- sp_relative_shift[uxn_opcodes_h_l1234_c30_ed5a] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_ins;
     sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_x;
     sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_return_output := sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1237_c21_c1f1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1237_c21_c1f1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c21_c1f1_left;
     BIN_OP_EQ_uxn_opcodes_h_l1237_c21_c1f1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c21_c1f1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c21_c1f1_return_output := BIN_OP_EQ_uxn_opcodes_h_l1237_c21_c1f1_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1218_c6_7b8d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1228_l1231_DUPLICATE_b093 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1228_l1231_DUPLICATE_b093_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1218_l1225_l1228_l1239_DUPLICATE_1934 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1218_l1225_l1228_l1239_DUPLICATE_1934_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1228_c11_fcc6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_left;
     BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_return_output := BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1218_l1225_l1228_l1239_DUPLICATE_bbcd LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1218_l1225_l1228_l1239_DUPLICATE_bbcd_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1239_c11_624d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1239_c11_624d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_624d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1239_c11_624d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_624d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_624d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1239_c11_624d_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1218_l1225_l1228_l1231_DUPLICATE_2373 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1218_l1225_l1228_l1231_DUPLICATE_2373_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1231_c11_8493] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493_left;
     BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493_return_output := BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1218_c2_4baf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1218_c2_4baf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1218_c6_7b8d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1225_c7_477a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1225_c7_477a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1225_c11_2770_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1228_c11_fcc6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c11_8493_return_output;
     VAR_MUX_uxn_opcodes_h_l1237_c21_e026_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1237_c21_c1f1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_624d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_624d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_624d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1218_l1225_l1228_l1239_DUPLICATE_1934_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1218_l1225_l1228_l1239_DUPLICATE_1934_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1218_l1225_l1228_l1239_DUPLICATE_1934_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1218_l1225_l1228_l1239_DUPLICATE_1934_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1239_l1225_l1228_l1231_DUPLICATE_0679_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1239_l1225_l1228_l1231_DUPLICATE_0679_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1239_l1225_l1228_l1231_DUPLICATE_0679_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1239_l1225_l1228_l1231_DUPLICATE_0679_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1218_l1225_l1228_l1239_DUPLICATE_bbcd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1218_l1225_l1228_l1239_DUPLICATE_bbcd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1218_l1225_l1228_l1239_DUPLICATE_bbcd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1218_l1225_l1228_l1239_DUPLICATE_bbcd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1228_l1231_DUPLICATE_b093_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1228_l1231_DUPLICATE_b093_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1218_l1225_l1228_l1231_DUPLICATE_2373_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1218_l1225_l1228_l1231_DUPLICATE_2373_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1218_l1225_l1228_l1231_DUPLICATE_2373_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1218_l1225_l1228_l1231_DUPLICATE_2373_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1234_c30_ed5a_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1239_c7_ddaa] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1239_c7_ddaa] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_return_output;

     -- MUX[uxn_opcodes_h_l1237_c21_e026] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1237_c21_e026_cond <= VAR_MUX_uxn_opcodes_h_l1237_c21_e026_cond;
     MUX_uxn_opcodes_h_l1237_c21_e026_iftrue <= VAR_MUX_uxn_opcodes_h_l1237_c21_e026_iftrue;
     MUX_uxn_opcodes_h_l1237_c21_e026_iffalse <= VAR_MUX_uxn_opcodes_h_l1237_c21_e026_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1237_c21_e026_return_output := MUX_uxn_opcodes_h_l1237_c21_e026_return_output;

     -- t8_MUX[uxn_opcodes_h_l1228_c7_ac0c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond <= VAR_t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond;
     t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue;
     t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output := t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1239_c7_ddaa] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1231_c7_5bf9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output;

     -- n8_MUX[uxn_opcodes_h_l1231_c7_5bf9] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond <= VAR_n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond;
     n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue;
     n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output := n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue := VAR_MUX_uxn_opcodes_h_l1237_c21_e026_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ddaa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ddaa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ddaa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output;
     -- t8_MUX[uxn_opcodes_h_l1225_c7_477a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1225_c7_477a_cond <= VAR_t8_MUX_uxn_opcodes_h_l1225_c7_477a_cond;
     t8_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue;
     t8_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1225_c7_477a_return_output := t8_MUX_uxn_opcodes_h_l1225_c7_477a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1228_c7_ac0c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output;

     -- n8_MUX[uxn_opcodes_h_l1228_c7_ac0c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond <= VAR_n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond;
     n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue;
     n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output := n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1231_c7_5bf9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1231_c7_5bf9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1231_c7_5bf9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1231_c7_5bf9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output := result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c7_5bf9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1225_c7_477a_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1228_c7_ac0c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1228_c7_ac0c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output;

     -- t8_MUX[uxn_opcodes_h_l1218_c2_4baf] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1218_c2_4baf_cond <= VAR_t8_MUX_uxn_opcodes_h_l1218_c2_4baf_cond;
     t8_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue;
     t8_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output := t8_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output;

     -- n8_MUX[uxn_opcodes_h_l1225_c7_477a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1225_c7_477a_cond <= VAR_n8_MUX_uxn_opcodes_h_l1225_c7_477a_cond;
     n8_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue;
     n8_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1225_c7_477a_return_output := n8_MUX_uxn_opcodes_h_l1225_c7_477a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1228_c7_ac0c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1225_c7_477a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1228_c7_ac0c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1225_c7_477a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1225_c7_477a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1228_c7_ac0c_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1225_c7_477a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1218_c2_4baf] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output;

     -- n8_MUX[uxn_opcodes_h_l1218_c2_4baf] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1218_c2_4baf_cond <= VAR_n8_MUX_uxn_opcodes_h_l1218_c2_4baf_cond;
     n8_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue;
     n8_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output := n8_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1225_c7_477a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1225_c7_477a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1225_c7_477a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_return_output := result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1225_c7_477a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1225_c7_477a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1225_c7_477a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1225_c7_477a_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1218_c2_4baf] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1218_c2_4baf] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1218_c2_4baf] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output := result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1218_c2_4baf] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1214_l1245_DUPLICATE_ab89 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1214_l1245_DUPLICATE_ab89_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_eae7(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1218_c2_4baf_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1214_l1245_DUPLICATE_ab89_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1214_l1245_DUPLICATE_ab89_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
