-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 50
entity jmp2_0CLK_8b7cd1f2 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jmp2_0CLK_8b7cd1f2;
architecture arch of jmp2_0CLK_8b7cd1f2 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l656_c6_3781]
signal BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l656_c2_c7b4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output : signed(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l656_c2_c7b4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output : unsigned(7 downto 0);

-- result_pc_MUX[uxn_opcodes_h_l656_c2_c7b4]
signal result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_cond : unsigned(0 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l656_c2_c7b4]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l656_c2_c7b4]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l656_c2_c7b4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l656_c2_c7b4]
signal t16_MUX_uxn_opcodes_h_l656_c2_c7b4_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l661_c11_342d]
signal BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l661_c7_5ea5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output : signed(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l661_c7_5ea5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output : unsigned(7 downto 0);

-- result_pc_MUX[uxn_opcodes_h_l661_c7_5ea5]
signal result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_cond : unsigned(0 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l661_c7_5ea5]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l661_c7_5ea5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l661_c7_5ea5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l661_c7_5ea5]
signal t16_MUX_uxn_opcodes_h_l661_c7_5ea5_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l664_c11_c4a8]
signal BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l664_c7_1754]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_return_output : signed(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l664_c7_1754]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_return_output : unsigned(7 downto 0);

-- result_pc_MUX[uxn_opcodes_h_l664_c7_1754]
signal result_pc_MUX_uxn_opcodes_h_l664_c7_1754_cond : unsigned(0 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l664_c7_1754_iftrue : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l664_c7_1754_iffalse : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l664_c7_1754_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l664_c7_1754]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l664_c7_1754]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l664_c7_1754]
signal result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l664_c7_1754]
signal t16_MUX_uxn_opcodes_h_l664_c7_1754_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l664_c7_1754_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l664_c7_1754_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l664_c7_1754_return_output : unsigned(15 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l666_c3_6f15]
signal CONST_SL_8_uxn_opcodes_h_l666_c3_6f15_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l666_c3_6f15_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l669_c11_97cc]
signal BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l669_c7_b0bd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output : signed(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l669_c7_b0bd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output : unsigned(7 downto 0);

-- result_pc_MUX[uxn_opcodes_h_l669_c7_b0bd]
signal result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_cond : unsigned(0 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l669_c7_b0bd]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l669_c7_b0bd]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l669_c7_b0bd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l669_c7_b0bd]
signal t16_MUX_uxn_opcodes_h_l669_c7_b0bd_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l672_c11_2b56]
signal BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l672_c7_2672]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_return_output : signed(7 downto 0);

-- result_pc_MUX[uxn_opcodes_h_l672_c7_2672]
signal result_pc_MUX_uxn_opcodes_h_l672_c7_2672_cond : unsigned(0 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l672_c7_2672_iftrue : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l672_c7_2672_iffalse : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l672_c7_2672_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l672_c7_2672]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l672_c7_2672]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l672_c7_2672]
signal result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l672_c7_2672]
signal t16_MUX_uxn_opcodes_h_l672_c7_2672_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l672_c7_2672_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l672_c7_2672_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l672_c7_2672_return_output : unsigned(15 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l673_c3_002e]
signal BIN_OP_OR_uxn_opcodes_h_l673_c3_002e_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l673_c3_002e_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l673_c3_002e_return_output : unsigned(15 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l675_c32_2476]
signal BIN_OP_AND_uxn_opcodes_h_l675_c32_2476_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l675_c32_2476_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l675_c32_2476_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l675_c32_cea4]
signal BIN_OP_GT_uxn_opcodes_h_l675_c32_cea4_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l675_c32_cea4_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l675_c32_cea4_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l675_c32_e328]
signal MUX_uxn_opcodes_h_l675_c32_e328_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l675_c32_e328_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l675_c32_e328_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l675_c32_e328_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l679_c11_0d1e]
signal BIN_OP_EQ_uxn_opcodes_h_l679_c11_0d1e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l679_c11_0d1e_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l679_c11_0d1e_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l679_c7_c67b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l679_c7_c67b]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l679_c7_c67b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_return_output : unsigned(0 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_f07d( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.pc := ref_toks_3;
      base.is_pc_updated := ref_toks_4;
      base.is_sp_shift := ref_toks_5;
      base.is_opc_done := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781
BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_left,
BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_right,
BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4
result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output);

-- result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4
result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_cond,
result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue,
result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse,
result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4
result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4
result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4
result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output);

-- t16_MUX_uxn_opcodes_h_l656_c2_c7b4
t16_MUX_uxn_opcodes_h_l656_c2_c7b4 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l656_c2_c7b4_cond,
t16_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue,
t16_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse,
t16_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d
BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_left,
BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_right,
BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5
result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output);

-- result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5
result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_cond,
result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue,
result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse,
result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5
result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5
result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5
result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output);

-- t16_MUX_uxn_opcodes_h_l661_c7_5ea5
t16_MUX_uxn_opcodes_h_l661_c7_5ea5 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l661_c7_5ea5_cond,
t16_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue,
t16_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse,
t16_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8
BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_left,
BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_right,
BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754
result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_return_output);

-- result_pc_MUX_uxn_opcodes_h_l664_c7_1754
result_pc_MUX_uxn_opcodes_h_l664_c7_1754 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_pc_MUX_uxn_opcodes_h_l664_c7_1754_cond,
result_pc_MUX_uxn_opcodes_h_l664_c7_1754_iftrue,
result_pc_MUX_uxn_opcodes_h_l664_c7_1754_iffalse,
result_pc_MUX_uxn_opcodes_h_l664_c7_1754_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754
result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754
result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754
result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_return_output);

-- t16_MUX_uxn_opcodes_h_l664_c7_1754
t16_MUX_uxn_opcodes_h_l664_c7_1754 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l664_c7_1754_cond,
t16_MUX_uxn_opcodes_h_l664_c7_1754_iftrue,
t16_MUX_uxn_opcodes_h_l664_c7_1754_iffalse,
t16_MUX_uxn_opcodes_h_l664_c7_1754_return_output);

-- CONST_SL_8_uxn_opcodes_h_l666_c3_6f15
CONST_SL_8_uxn_opcodes_h_l666_c3_6f15 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l666_c3_6f15_x,
CONST_SL_8_uxn_opcodes_h_l666_c3_6f15_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc
BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_left,
BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_right,
BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd
result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output);

-- result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd
result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_cond,
result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue,
result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse,
result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd
result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd
result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd
result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output);

-- t16_MUX_uxn_opcodes_h_l669_c7_b0bd
t16_MUX_uxn_opcodes_h_l669_c7_b0bd : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l669_c7_b0bd_cond,
t16_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue,
t16_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse,
t16_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56
BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56_left,
BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56_right,
BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672
result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_return_output);

-- result_pc_MUX_uxn_opcodes_h_l672_c7_2672
result_pc_MUX_uxn_opcodes_h_l672_c7_2672 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_pc_MUX_uxn_opcodes_h_l672_c7_2672_cond,
result_pc_MUX_uxn_opcodes_h_l672_c7_2672_iftrue,
result_pc_MUX_uxn_opcodes_h_l672_c7_2672_iffalse,
result_pc_MUX_uxn_opcodes_h_l672_c7_2672_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672
result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672
result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672
result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_return_output);

-- t16_MUX_uxn_opcodes_h_l672_c7_2672
t16_MUX_uxn_opcodes_h_l672_c7_2672 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l672_c7_2672_cond,
t16_MUX_uxn_opcodes_h_l672_c7_2672_iftrue,
t16_MUX_uxn_opcodes_h_l672_c7_2672_iffalse,
t16_MUX_uxn_opcodes_h_l672_c7_2672_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l673_c3_002e
BIN_OP_OR_uxn_opcodes_h_l673_c3_002e : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l673_c3_002e_left,
BIN_OP_OR_uxn_opcodes_h_l673_c3_002e_right,
BIN_OP_OR_uxn_opcodes_h_l673_c3_002e_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l675_c32_2476
BIN_OP_AND_uxn_opcodes_h_l675_c32_2476 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l675_c32_2476_left,
BIN_OP_AND_uxn_opcodes_h_l675_c32_2476_right,
BIN_OP_AND_uxn_opcodes_h_l675_c32_2476_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l675_c32_cea4
BIN_OP_GT_uxn_opcodes_h_l675_c32_cea4 : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l675_c32_cea4_left,
BIN_OP_GT_uxn_opcodes_h_l675_c32_cea4_right,
BIN_OP_GT_uxn_opcodes_h_l675_c32_cea4_return_output);

-- MUX_uxn_opcodes_h_l675_c32_e328
MUX_uxn_opcodes_h_l675_c32_e328 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l675_c32_e328_cond,
MUX_uxn_opcodes_h_l675_c32_e328_iftrue,
MUX_uxn_opcodes_h_l675_c32_e328_iffalse,
MUX_uxn_opcodes_h_l675_c32_e328_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l679_c11_0d1e
BIN_OP_EQ_uxn_opcodes_h_l679_c11_0d1e : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l679_c11_0d1e_left,
BIN_OP_EQ_uxn_opcodes_h_l679_c11_0d1e_right,
BIN_OP_EQ_uxn_opcodes_h_l679_c11_0d1e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b
result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b
result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b
result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output,
 result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output,
 t16_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output,
 result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output,
 t16_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_return_output,
 result_pc_MUX_uxn_opcodes_h_l664_c7_1754_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_return_output,
 t16_MUX_uxn_opcodes_h_l664_c7_1754_return_output,
 CONST_SL_8_uxn_opcodes_h_l666_c3_6f15_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output,
 result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output,
 t16_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_return_output,
 result_pc_MUX_uxn_opcodes_h_l672_c7_2672_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_return_output,
 t16_MUX_uxn_opcodes_h_l672_c7_2672_return_output,
 BIN_OP_OR_uxn_opcodes_h_l673_c3_002e_return_output,
 BIN_OP_AND_uxn_opcodes_h_l675_c32_2476_return_output,
 BIN_OP_GT_uxn_opcodes_h_l675_c32_cea4_return_output,
 MUX_uxn_opcodes_h_l675_c32_e328_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l679_c11_0d1e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l658_c3_1b41 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_cond : unsigned(0 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l656_c2_c7b4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l662_c3_2cbf : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_cond : unsigned(0 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l664_c7_1754_return_output : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l664_c7_1754_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l661_c7_5ea5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l667_c3_5338 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_cond : unsigned(0 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l664_c7_1754_iftrue : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l664_c7_1754_iffalse : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l664_c7_1754_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l664_c7_1754_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l664_c7_1754_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l664_c7_1754_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l666_c3_6f15_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l666_c3_6f15_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l670_c3_9db9 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l669_c7_b0bd_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_cond : unsigned(0 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l672_c7_2672_return_output : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l672_c7_2672_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l669_c7_b0bd_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_cond : unsigned(0 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l672_c7_2672_iftrue : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l672_c7_2672_iffalse : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l672_c7_2672_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l672_c7_2672_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l672_c7_2672_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l672_c7_2672_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l673_c3_002e_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l673_c3_002e_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l673_c3_002e_return_output : unsigned(15 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l675_c32_e328_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l675_c32_e328_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l675_c32_e328_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l675_c32_2476_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l675_c32_2476_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l675_c32_2476_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l675_c32_cea4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l675_c32_cea4_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l675_c32_cea4_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l675_c32_e328_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l679_c11_0d1e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l679_c11_0d1e_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l679_c11_0d1e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l661_l672_l656_l669_l664_DUPLICATE_e367_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l661_l672_l656_l669_l664_DUPLICATE_fecd_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l661_l679_l656_l669_l664_DUPLICATE_028f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l661_l679_l656_l669_l664_DUPLICATE_cd0b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l661_l679_l672_l669_l664_DUPLICATE_ea93_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l665_l673_DUPLICATE_ce9d_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_f07d_uxn_opcodes_h_l652_l685_DUPLICATE_5f43_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l679_c11_0d1e_right := to_unsigned(5, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l658_c3_1b41 := resize(to_unsigned(2, 2), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l658_c3_1b41;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l667_c3_5338 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l667_c3_5338;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l670_c3_9db9 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l670_c3_9db9;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l662_c3_2cbf := resize(to_unsigned(2, 2), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l662_c3_2cbf;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_right := to_unsigned(3, 2);
     VAR_BIN_OP_AND_uxn_opcodes_h_l675_c32_2476_right := to_unsigned(128, 8);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_right := to_unsigned(0, 1);
     VAR_BIN_OP_GT_uxn_opcodes_h_l675_c32_cea4_right := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l675_c32_e328_iftrue := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_MUX_uxn_opcodes_h_l675_c32_e328_iffalse := resize(to_signed(-2, 3), 8);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_BIN_OP_AND_uxn_opcodes_h_l675_c32_2476_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l679_c11_0d1e_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l673_c3_002e_left := t16;
     VAR_t16_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l672_c7_2672_iffalse := t16;
     -- BIN_OP_EQ[uxn_opcodes_h_l664_c11_c4a8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_left;
     BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_return_output := BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_return_output;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l661_l672_l656_l669_l664_DUPLICATE_e367 LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l661_l672_l656_l669_l664_DUPLICATE_e367_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l661_l672_l656_l669_l664_DUPLICATE_fecd LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l661_l672_l656_l669_l664_DUPLICATE_fecd_return_output := result.pc;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l661_l679_l656_l669_l664_DUPLICATE_cd0b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l661_l679_l656_l669_l664_DUPLICATE_cd0b_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l679_c11_0d1e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l679_c11_0d1e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l679_c11_0d1e_left;
     BIN_OP_EQ_uxn_opcodes_h_l679_c11_0d1e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l679_c11_0d1e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l679_c11_0d1e_return_output := BIN_OP_EQ_uxn_opcodes_h_l679_c11_0d1e_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l669_c7_b0bd] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l669_c7_b0bd_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l672_c11_2b56] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56_left;
     BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56_return_output := BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l661_l679_l656_l669_l664_DUPLICATE_028f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l661_l679_l656_l669_l664_DUPLICATE_028f_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l669_c11_97cc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_left;
     BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_return_output := BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l661_l679_l672_l669_l664_DUPLICATE_ea93 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l661_l679_l672_l669_l664_DUPLICATE_ea93_return_output := result.is_opc_done;

     -- BIN_OP_AND[uxn_opcodes_h_l675_c32_2476] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l675_c32_2476_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l675_c32_2476_left;
     BIN_OP_AND_uxn_opcodes_h_l675_c32_2476_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l675_c32_2476_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l675_c32_2476_return_output := BIN_OP_AND_uxn_opcodes_h_l675_c32_2476_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l661_c11_342d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_left;
     BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_return_output := BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_return_output;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l665_l673_DUPLICATE_ce9d LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l665_l673_DUPLICATE_ce9d_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l656_c6_3781] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_left;
     BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_return_output := BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_return_output;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l675_c32_cea4_left := VAR_BIN_OP_AND_uxn_opcodes_h_l675_c32_2476_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l656_c2_c7b4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_3781_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l661_c7_5ea5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_342d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l664_c7_1754_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l664_c7_1754_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_c4a8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l669_c7_b0bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_97cc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l672_c7_2672_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l672_c7_2672_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_2b56_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l679_c11_0d1e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l679_c11_0d1e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l679_c11_0d1e_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l673_c3_002e_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l665_l673_DUPLICATE_ce9d_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l666_c3_6f15_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l665_l673_DUPLICATE_ce9d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l661_l672_l656_l669_l664_DUPLICATE_e367_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l661_l672_l656_l669_l664_DUPLICATE_e367_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l661_l672_l656_l669_l664_DUPLICATE_e367_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l661_l672_l656_l669_l664_DUPLICATE_e367_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l661_l672_l656_l669_l664_DUPLICATE_e367_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l661_l672_l656_l669_l664_DUPLICATE_fecd_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l661_l672_l656_l669_l664_DUPLICATE_fecd_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l664_c7_1754_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l661_l672_l656_l669_l664_DUPLICATE_fecd_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l661_l672_l656_l669_l664_DUPLICATE_fecd_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l672_c7_2672_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l661_l672_l656_l669_l664_DUPLICATE_fecd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l661_l679_l672_l669_l664_DUPLICATE_ea93_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l661_l679_l672_l669_l664_DUPLICATE_ea93_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l661_l679_l672_l669_l664_DUPLICATE_ea93_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l661_l679_l672_l669_l664_DUPLICATE_ea93_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l661_l679_l672_l669_l664_DUPLICATE_ea93_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l661_l679_l656_l669_l664_DUPLICATE_028f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l661_l679_l656_l669_l664_DUPLICATE_028f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l661_l679_l656_l669_l664_DUPLICATE_028f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l661_l679_l656_l669_l664_DUPLICATE_028f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l661_l679_l656_l669_l664_DUPLICATE_028f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l661_l679_l656_l669_l664_DUPLICATE_cd0b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l661_l679_l656_l669_l664_DUPLICATE_cd0b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l661_l679_l656_l669_l664_DUPLICATE_cd0b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l661_l679_l656_l669_l664_DUPLICATE_cd0b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l661_l679_l656_l669_l664_DUPLICATE_cd0b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l669_c7_b0bd_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l669_c7_b0bd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l673_c3_002e] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l673_c3_002e_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l673_c3_002e_left;
     BIN_OP_OR_uxn_opcodes_h_l673_c3_002e_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l673_c3_002e_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l673_c3_002e_return_output := BIN_OP_OR_uxn_opcodes_h_l673_c3_002e_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l666_c3_6f15] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l666_c3_6f15_x <= VAR_CONST_SL_8_uxn_opcodes_h_l666_c3_6f15_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l666_c3_6f15_return_output := CONST_SL_8_uxn_opcodes_h_l666_c3_6f15_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l679_c7_c67b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l679_c7_c67b] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l675_c32_cea4] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l675_c32_cea4_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l675_c32_cea4_left;
     BIN_OP_GT_uxn_opcodes_h_l675_c32_cea4_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l675_c32_cea4_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l675_c32_cea4_return_output := BIN_OP_GT_uxn_opcodes_h_l675_c32_cea4_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l679_c7_c67b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l675_c32_e328_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l675_c32_cea4_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l672_c7_2672_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l673_c3_002e_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l672_c7_2672_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l673_c3_002e_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l664_c7_1754_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l666_c3_6f15_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_c67b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_c67b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_c67b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output;
     -- result_pc_MUX[uxn_opcodes_h_l672_c7_2672] LATENCY=0
     -- Inputs
     result_pc_MUX_uxn_opcodes_h_l672_c7_2672_cond <= VAR_result_pc_MUX_uxn_opcodes_h_l672_c7_2672_cond;
     result_pc_MUX_uxn_opcodes_h_l672_c7_2672_iftrue <= VAR_result_pc_MUX_uxn_opcodes_h_l672_c7_2672_iftrue;
     result_pc_MUX_uxn_opcodes_h_l672_c7_2672_iffalse <= VAR_result_pc_MUX_uxn_opcodes_h_l672_c7_2672_iffalse;
     -- Outputs
     VAR_result_pc_MUX_uxn_opcodes_h_l672_c7_2672_return_output := result_pc_MUX_uxn_opcodes_h_l672_c7_2672_return_output;

     -- MUX[uxn_opcodes_h_l675_c32_e328] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l675_c32_e328_cond <= VAR_MUX_uxn_opcodes_h_l675_c32_e328_cond;
     MUX_uxn_opcodes_h_l675_c32_e328_iftrue <= VAR_MUX_uxn_opcodes_h_l675_c32_e328_iftrue;
     MUX_uxn_opcodes_h_l675_c32_e328_iffalse <= VAR_MUX_uxn_opcodes_h_l675_c32_e328_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l675_c32_e328_return_output := MUX_uxn_opcodes_h_l675_c32_e328_return_output;

     -- t16_MUX[uxn_opcodes_h_l672_c7_2672] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l672_c7_2672_cond <= VAR_t16_MUX_uxn_opcodes_h_l672_c7_2672_cond;
     t16_MUX_uxn_opcodes_h_l672_c7_2672_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l672_c7_2672_iftrue;
     t16_MUX_uxn_opcodes_h_l672_c7_2672_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l672_c7_2672_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l672_c7_2672_return_output := t16_MUX_uxn_opcodes_h_l672_c7_2672_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l664_c7_1754] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l672_c7_2672] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l672_c7_2672] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l672_c7_2672] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_iftrue := VAR_MUX_uxn_opcodes_h_l675_c32_e328_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_2672_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_2672_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_2672_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse := VAR_result_pc_MUX_uxn_opcodes_h_l672_c7_2672_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_1754_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse := VAR_t16_MUX_uxn_opcodes_h_l672_c7_2672_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l669_c7_b0bd] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output;

     -- result_pc_MUX[uxn_opcodes_h_l669_c7_b0bd] LATENCY=0
     -- Inputs
     result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_cond <= VAR_result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_cond;
     result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue <= VAR_result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue;
     result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse <= VAR_result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse;
     -- Outputs
     VAR_result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output := result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l669_c7_b0bd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l672_c7_2672] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l669_c7_b0bd] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output;

     -- t16_MUX[uxn_opcodes_h_l669_c7_b0bd] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l669_c7_b0bd_cond <= VAR_t16_MUX_uxn_opcodes_h_l669_c7_b0bd_cond;
     t16_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue;
     t16_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output := t16_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l661_c7_5ea5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l664_c7_1754_iffalse := VAR_result_pc_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_2672_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l664_c7_1754_iffalse := VAR_t16_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l664_c7_1754] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_return_output;

     -- result_pc_MUX[uxn_opcodes_h_l664_c7_1754] LATENCY=0
     -- Inputs
     result_pc_MUX_uxn_opcodes_h_l664_c7_1754_cond <= VAR_result_pc_MUX_uxn_opcodes_h_l664_c7_1754_cond;
     result_pc_MUX_uxn_opcodes_h_l664_c7_1754_iftrue <= VAR_result_pc_MUX_uxn_opcodes_h_l664_c7_1754_iftrue;
     result_pc_MUX_uxn_opcodes_h_l664_c7_1754_iffalse <= VAR_result_pc_MUX_uxn_opcodes_h_l664_c7_1754_iffalse;
     -- Outputs
     VAR_result_pc_MUX_uxn_opcodes_h_l664_c7_1754_return_output := result_pc_MUX_uxn_opcodes_h_l664_c7_1754_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l664_c7_1754] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l656_c2_c7b4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output;

     -- t16_MUX[uxn_opcodes_h_l664_c7_1754] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l664_c7_1754_cond <= VAR_t16_MUX_uxn_opcodes_h_l664_c7_1754_cond;
     t16_MUX_uxn_opcodes_h_l664_c7_1754_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l664_c7_1754_iftrue;
     t16_MUX_uxn_opcodes_h_l664_c7_1754_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l664_c7_1754_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l664_c7_1754_return_output := t16_MUX_uxn_opcodes_h_l664_c7_1754_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l669_c7_b0bd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l664_c7_1754] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_1754_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_1754_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_1754_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse := VAR_result_pc_MUX_uxn_opcodes_h_l664_c7_1754_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_b0bd_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse := VAR_t16_MUX_uxn_opcodes_h_l664_c7_1754_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l661_c7_5ea5] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l661_c7_5ea5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l664_c7_1754] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_return_output;

     -- result_pc_MUX[uxn_opcodes_h_l661_c7_5ea5] LATENCY=0
     -- Inputs
     result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_cond <= VAR_result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_cond;
     result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue <= VAR_result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue;
     result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse <= VAR_result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse;
     -- Outputs
     VAR_result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output := result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l661_c7_5ea5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output;

     -- t16_MUX[uxn_opcodes_h_l661_c7_5ea5] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l661_c7_5ea5_cond <= VAR_t16_MUX_uxn_opcodes_h_l661_c7_5ea5_cond;
     t16_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue;
     t16_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output := t16_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse := VAR_result_pc_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_1754_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse := VAR_t16_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output;
     -- result_pc_MUX[uxn_opcodes_h_l656_c2_c7b4] LATENCY=0
     -- Inputs
     result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_cond <= VAR_result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_cond;
     result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue <= VAR_result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue;
     result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse <= VAR_result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse;
     -- Outputs
     VAR_result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output := result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l656_c2_c7b4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l656_c2_c7b4] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output;

     -- t16_MUX[uxn_opcodes_h_l656_c2_c7b4] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l656_c2_c7b4_cond <= VAR_t16_MUX_uxn_opcodes_h_l656_c2_c7b4_cond;
     t16_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue;
     t16_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output := t16_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l656_c2_c7b4] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l661_c7_5ea5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output;

     -- Submodule level 7
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_5ea5_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l656_c2_c7b4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output;

     -- Submodule level 8
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_f07d_uxn_opcodes_h_l652_l685_DUPLICATE_5f43 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_f07d_uxn_opcodes_h_l652_l685_DUPLICATE_5f43_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_f07d(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output,
     VAR_result_pc_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_c7b4_return_output);

     -- Submodule level 9
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_f07d_uxn_opcodes_h_l652_l685_DUPLICATE_5f43_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_f07d_uxn_opcodes_h_l652_l685_DUPLICATE_5f43_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
