-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 55
entity lit2_0CLK_edc09f97 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end lit2_0CLK_edc09f97;
architecture arch of lit2_0CLK_edc09f97 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal tmp16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_tmp16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l214_c6_074e]
signal BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l214_c1_2c16]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l214_c2_9f76]
signal tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l214_c2_9f76]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l214_c2_9f76]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l214_c2_9f76]
signal result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l214_c2_9f76]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l214_c2_9f76]
signal result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l214_c2_9f76]
signal result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_return_output : unsigned(15 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l214_c2_9f76]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l214_c2_9f76]
signal result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l215_c3_6650[uxn_opcodes_h_l215_c3_6650]
signal printf_uxn_opcodes_h_l215_c3_6650_uxn_opcodes_h_l215_c3_6650_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l221_c11_1e7e]
signal BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l221_c7_3793]
signal tmp16_MUX_uxn_opcodes_h_l221_c7_3793_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l221_c7_3793_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l221_c7_3793_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l221_c7_3793_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l221_c7_3793]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l221_c7_3793]
signal result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l221_c7_3793]
signal result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l221_c7_3793]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l221_c7_3793]
signal result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l221_c7_3793]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l221_c7_3793]
signal result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_return_output : unsigned(7 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l223_c22_c5a0]
signal BIN_OP_PLUS_uxn_opcodes_h_l223_c22_c5a0_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l223_c22_c5a0_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l223_c22_c5a0_return_output : unsigned(16 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l225_c11_5454]
signal BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l225_c7_b145]
signal tmp16_MUX_uxn_opcodes_h_l225_c7_b145_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l225_c7_b145_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l225_c7_b145_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l225_c7_b145_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l225_c7_b145]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l225_c7_b145]
signal result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l225_c7_b145]
signal result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l225_c7_b145]
signal result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l225_c7_b145]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l225_c7_b145]
signal result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_return_output : unsigned(7 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l227_c3_14a4]
signal CONST_SL_8_uxn_opcodes_h_l227_c3_14a4_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l227_c3_14a4_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l229_c11_dffc]
signal BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l229_c7_ca0b]
signal tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l229_c7_ca0b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l229_c7_ca0b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l229_c7_ca0b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l229_c7_ca0b]
signal result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l229_c7_ca0b]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l229_c7_ca0b]
signal result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output : unsigned(7 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l230_c3_0c06]
signal BIN_OP_OR_uxn_opcodes_h_l230_c3_0c06_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l230_c3_0c06_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l230_c3_0c06_return_output : unsigned(15 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l232_c22_1ba2]
signal BIN_OP_PLUS_uxn_opcodes_h_l232_c22_1ba2_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l232_c22_1ba2_right : unsigned(1 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l232_c22_1ba2_return_output : unsigned(16 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l237_c11_0129]
signal BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l237_c7_7773]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l237_c7_7773]
signal result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l237_c7_7773]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l237_c7_7773]
signal result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l237_c7_7773]
signal result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_return_output : unsigned(7 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l240_c31_da49]
signal CONST_SR_8_uxn_opcodes_h_l240_c31_da49_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l240_c31_da49_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l242_c11_6c49]
signal BIN_OP_EQ_uxn_opcodes_h_l242_c11_6c49_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l242_c11_6c49_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l242_c11_6c49_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l242_c7_387e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l242_c7_387e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_return_output : unsigned(0 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_e2b8( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : signed;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.sp_relative_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_pc_updated := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.u16_value := ref_toks_6;
      base.is_sp_shift := ref_toks_7;
      base.u8_value := ref_toks_8;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e
BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_left,
BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_right,
BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_return_output);

-- tmp16_MUX_uxn_opcodes_h_l214_c2_9f76
tmp16_MUX_uxn_opcodes_h_l214_c2_9f76 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_cond,
tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue,
tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse,
tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76
result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76
result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76
result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76
result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76
result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_cond,
result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76
result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76
result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_cond,
result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_return_output);

-- printf_uxn_opcodes_h_l215_c3_6650_uxn_opcodes_h_l215_c3_6650
printf_uxn_opcodes_h_l215_c3_6650_uxn_opcodes_h_l215_c3_6650 : entity work.printf_uxn_opcodes_h_l215_c3_6650_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l215_c3_6650_uxn_opcodes_h_l215_c3_6650_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e
BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_left,
BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_right,
BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_return_output);

-- tmp16_MUX_uxn_opcodes_h_l221_c7_3793
tmp16_MUX_uxn_opcodes_h_l221_c7_3793 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l221_c7_3793_cond,
tmp16_MUX_uxn_opcodes_h_l221_c7_3793_iftrue,
tmp16_MUX_uxn_opcodes_h_l221_c7_3793_iffalse,
tmp16_MUX_uxn_opcodes_h_l221_c7_3793_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793
result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793
result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793
result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793
result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_cond,
result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793
result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793
result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_cond,
result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l223_c22_c5a0
BIN_OP_PLUS_uxn_opcodes_h_l223_c22_c5a0 : entity work.BIN_OP_PLUS_uint16_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l223_c22_c5a0_left,
BIN_OP_PLUS_uxn_opcodes_h_l223_c22_c5a0_right,
BIN_OP_PLUS_uxn_opcodes_h_l223_c22_c5a0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454
BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_left,
BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_right,
BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_return_output);

-- tmp16_MUX_uxn_opcodes_h_l225_c7_b145
tmp16_MUX_uxn_opcodes_h_l225_c7_b145 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l225_c7_b145_cond,
tmp16_MUX_uxn_opcodes_h_l225_c7_b145_iftrue,
tmp16_MUX_uxn_opcodes_h_l225_c7_b145_iffalse,
tmp16_MUX_uxn_opcodes_h_l225_c7_b145_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145
result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145
result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145
result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_cond,
result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145
result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145
result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_cond,
result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_return_output);

-- CONST_SL_8_uxn_opcodes_h_l227_c3_14a4
CONST_SL_8_uxn_opcodes_h_l227_c3_14a4 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l227_c3_14a4_x,
CONST_SL_8_uxn_opcodes_h_l227_c3_14a4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc
BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_left,
BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_right,
BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_return_output);

-- tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b
tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_cond,
tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue,
tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse,
tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b
result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b
result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b
result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_cond,
result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b
result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b
result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_cond,
result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l230_c3_0c06
BIN_OP_OR_uxn_opcodes_h_l230_c3_0c06 : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l230_c3_0c06_left,
BIN_OP_OR_uxn_opcodes_h_l230_c3_0c06_right,
BIN_OP_OR_uxn_opcodes_h_l230_c3_0c06_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l232_c22_1ba2
BIN_OP_PLUS_uxn_opcodes_h_l232_c22_1ba2 : entity work.BIN_OP_PLUS_uint16_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l232_c22_1ba2_left,
BIN_OP_PLUS_uxn_opcodes_h_l232_c22_1ba2_right,
BIN_OP_PLUS_uxn_opcodes_h_l232_c22_1ba2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129
BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129_left,
BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129_right,
BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773
result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773
result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773
result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773
result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_cond,
result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_return_output);

-- CONST_SR_8_uxn_opcodes_h_l240_c31_da49
CONST_SR_8_uxn_opcodes_h_l240_c31_da49 : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l240_c31_da49_x,
CONST_SR_8_uxn_opcodes_h_l240_c31_da49_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l242_c11_6c49
BIN_OP_EQ_uxn_opcodes_h_l242_c11_6c49 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l242_c11_6c49_left,
BIN_OP_EQ_uxn_opcodes_h_l242_c11_6c49_right,
BIN_OP_EQ_uxn_opcodes_h_l242_c11_6c49_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e
result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e
result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 previous_ram_read,
 -- Registers
 tmp16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_return_output,
 tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_return_output,
 tmp16_MUX_uxn_opcodes_h_l221_c7_3793_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l223_c22_c5a0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_return_output,
 tmp16_MUX_uxn_opcodes_h_l225_c7_b145_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_return_output,
 CONST_SL_8_uxn_opcodes_h_l227_c3_14a4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_return_output,
 tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output,
 BIN_OP_OR_uxn_opcodes_h_l230_c3_0c06_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l232_c22_1ba2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_return_output,
 CONST_SR_8_uxn_opcodes_h_l240_c31_da49_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l242_c11_6c49_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_iffalse : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_3793_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l217_c3_6706 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l214_c2_9f76_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l215_c3_6650_uxn_opcodes_h_l215_c3_6650_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_3793_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_3793_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_b145_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_3793_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l221_c7_3793_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l223_c3_8c5d : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_c5a0_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_c5a0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_c5a0_return_output : unsigned(16 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_b145_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_b145_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_b145_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l227_c3_14a4_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l227_c3_14a4_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l234_c3_5f0f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l232_c3_70b3 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_0c06_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_0c06_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_0c06_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_1ba2_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_1ba2_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_1ba2_return_output : unsigned(16 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l235_c21_f831_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l239_c3_fe01 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l240_c31_da49_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l240_c31_da49_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l240_c21_6b06_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_6c49_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_6c49_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_6c49_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l225_l214_l221_l237_DUPLICATE_a758_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l225_l214_l221_l237_DUPLICATE_40fb_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l225_l221_l214_l242_l237_DUPLICATE_ae10_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l225_l214_l221_l237_DUPLICATE_a609_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l225_l221_l242_l237_l229_DUPLICATE_f395_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l226_l230_DUPLICATE_d594_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l225_l229_DUPLICATE_07c4_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e2b8_uxn_opcodes_h_l247_l209_DUPLICATE_d25b_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_tmp16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_tmp16 := tmp16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_1ba2_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_right := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_iffalse := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_6c49_right := to_unsigned(5, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l239_c3_fe01 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l239_c3_fe01;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l217_c3_6706 := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l217_c3_6706;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l234_c3_5f0f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l234_c3_5f0f;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_c5a0_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_right := to_unsigned(3, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129_right := to_unsigned(4, 3);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_c5a0_left := VAR_pc;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_1ba2_left := VAR_pc;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_6c49_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_0c06_left := tmp16;
     VAR_CONST_SR_8_uxn_opcodes_h_l240_c31_da49_x := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_3793_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse := tmp16;
     -- BIN_OP_EQ[uxn_opcodes_h_l242_c11_6c49] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l242_c11_6c49_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_6c49_left;
     BIN_OP_EQ_uxn_opcodes_h_l242_c11_6c49_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_6c49_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_6c49_return_output := BIN_OP_EQ_uxn_opcodes_h_l242_c11_6c49_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l225_l214_l221_l237_DUPLICATE_a609 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l225_l214_l221_l237_DUPLICATE_a609_return_output := result.u8_value;

     -- result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d[uxn_opcodes_h_l214_c2_9f76] LATENCY=0
     VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l214_c2_9f76_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l237_c11_0129] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129_left;
     BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129_return_output := BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l229_c11_dffc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_left;
     BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_return_output := BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l225_l229_DUPLICATE_07c4 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l225_l229_DUPLICATE_07c4_return_output := result.u16_value;

     -- BIN_OP_PLUS[uxn_opcodes_h_l223_c22_c5a0] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l223_c22_c5a0_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_c5a0_left;
     BIN_OP_PLUS_uxn_opcodes_h_l223_c22_c5a0_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_c5a0_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_c5a0_return_output := BIN_OP_PLUS_uxn_opcodes_h_l223_c22_c5a0_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l225_l214_l221_l237_DUPLICATE_40fb LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l225_l214_l221_l237_DUPLICATE_40fb_return_output := result.is_pc_updated;

     -- BIN_OP_PLUS[uxn_opcodes_h_l232_c22_1ba2] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l232_c22_1ba2_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_1ba2_left;
     BIN_OP_PLUS_uxn_opcodes_h_l232_c22_1ba2_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_1ba2_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_1ba2_return_output := BIN_OP_PLUS_uxn_opcodes_h_l232_c22_1ba2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l225_c11_5454] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_left;
     BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_return_output := BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_return_output;

     -- result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d[uxn_opcodes_h_l221_c7_3793] LATENCY=0
     VAR_result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l221_c7_3793_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l221_c11_1e7e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_left;
     BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_return_output := BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l225_l221_l242_l237_l229_DUPLICATE_f395 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l225_l221_l242_l237_l229_DUPLICATE_f395_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l214_c6_074e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_left;
     BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_return_output := BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l225_l221_l214_l242_l237_DUPLICATE_ae10 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l225_l221_l214_l242_l237_DUPLICATE_ae10_return_output := result.is_stack_write;

     -- CONST_SR_8[uxn_opcodes_h_l240_c31_da49] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l240_c31_da49_x <= VAR_CONST_SR_8_uxn_opcodes_h_l240_c31_da49_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l240_c31_da49_return_output := CONST_SR_8_uxn_opcodes_h_l240_c31_da49_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l225_l214_l221_l237_DUPLICATE_a758 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l225_l214_l221_l237_DUPLICATE_a758_return_output := result.stack_address_sp_offset;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l226_l230_DUPLICATE_d594 LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l226_l230_DUPLICATE_d594_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_ram_read);

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_074e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_3793_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_1e7e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_b145_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_5454_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_dffc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_0129_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_6c49_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_6c49_return_output;
     VAR_result_u16_value_uxn_opcodes_h_l223_c3_8c5d := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_c5a0_return_output, 16);
     VAR_result_u16_value_uxn_opcodes_h_l232_c3_70b3 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_1ba2_return_output, 16);
     VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_0c06_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l226_l230_DUPLICATE_d594_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l227_c3_14a4_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l226_l230_DUPLICATE_d594_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l225_l229_DUPLICATE_07c4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l225_l229_DUPLICATE_07c4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l225_l221_l242_l237_l229_DUPLICATE_f395_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l225_l221_l242_l237_l229_DUPLICATE_f395_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l225_l221_l242_l237_l229_DUPLICATE_f395_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l225_l221_l242_l237_l229_DUPLICATE_f395_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l225_l221_l242_l237_l229_DUPLICATE_f395_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l225_l214_l221_l237_DUPLICATE_40fb_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l225_l214_l221_l237_DUPLICATE_40fb_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l225_l214_l221_l237_DUPLICATE_40fb_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l225_l214_l221_l237_DUPLICATE_40fb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l225_l221_l214_l242_l237_DUPLICATE_ae10_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l225_l221_l214_l242_l237_DUPLICATE_ae10_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l225_l221_l214_l242_l237_DUPLICATE_ae10_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l225_l221_l214_l242_l237_DUPLICATE_ae10_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l225_l221_l214_l242_l237_DUPLICATE_ae10_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l225_l214_l221_l237_DUPLICATE_a758_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l225_l214_l221_l237_DUPLICATE_a758_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l225_l214_l221_l237_DUPLICATE_a758_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l225_l214_l221_l237_DUPLICATE_a758_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l225_l214_l221_l237_DUPLICATE_a609_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l225_l214_l221_l237_DUPLICATE_a609_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l225_l214_l221_l237_DUPLICATE_a609_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l225_l214_l221_l237_DUPLICATE_a609_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_iffalse := VAR_result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l221_c7_3793_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse := VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l214_c2_9f76_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_iftrue := VAR_result_u16_value_uxn_opcodes_h_l223_c3_8c5d;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue := VAR_result_u16_value_uxn_opcodes_h_l232_c3_70b3;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l221_c7_3793] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l214_c2_9f76] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l214_c1_2c16] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l237_c7_7773] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l242_c7_387e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l229_c7_ca0b] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_cond;
     result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output := result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l230_c3_0c06] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l230_c3_0c06_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_0c06_left;
     BIN_OP_OR_uxn_opcodes_h_l230_c3_0c06_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_0c06_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_0c06_return_output := BIN_OP_OR_uxn_opcodes_h_l230_c3_0c06_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l242_c7_387e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l237_c7_7773] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l227_c3_14a4] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l227_c3_14a4_x <= VAR_CONST_SL_8_uxn_opcodes_h_l227_c3_14a4_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l227_c3_14a4_return_output := CONST_SL_8_uxn_opcodes_h_l227_c3_14a4_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l240_c21_6b06] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l240_c21_6b06_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l240_c31_da49_return_output);

     -- Submodule level 2
     VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_0c06_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l240_c21_6b06_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_b145_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l227_c3_14a4_return_output;
     VAR_printf_uxn_opcodes_h_l215_c3_6650_uxn_opcodes_h_l215_c3_6650_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_2c16_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_387e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_7773_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_3793_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_387e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_7773_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l214_c2_9f76] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l225_c7_b145] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_cond;
     result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_return_output := result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l229_c7_ca0b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l235_c21_f831] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l235_c21_f831_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_0c06_return_output);

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l229_c7_ca0b] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l237_c7_7773] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l237_c7_7773] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_cond;
     result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_return_output := result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l229_c7_ca0b] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_cond;
     tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue;
     tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output := tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l237_c7_7773] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_return_output;

     -- printf_uxn_opcodes_h_l215_c3_6650[uxn_opcodes_h_l215_c3_6650] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l215_c3_6650_uxn_opcodes_h_l215_c3_6650_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l215_c3_6650_uxn_opcodes_h_l215_c3_6650_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- Submodule level 3
     VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l235_c21_f831_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_7773_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_7773_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_b145_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_7773_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_b145_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l229_c7_ca0b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l229_c7_ca0b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l225_c7_b145] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l225_c7_b145_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_b145_cond;
     tmp16_MUX_uxn_opcodes_h_l225_c7_b145_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_b145_iftrue;
     tmp16_MUX_uxn_opcodes_h_l225_c7_b145_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_b145_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_b145_return_output := tmp16_MUX_uxn_opcodes_h_l225_c7_b145_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l225_c7_b145] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l229_c7_ca0b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output := result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l221_c7_3793] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_cond;
     result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_return_output := result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l225_c7_b145] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b145_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b145_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_3793_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_ca0b_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_3793_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_b145_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l225_c7_b145] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_cond;
     result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_return_output := result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l225_c7_b145] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l221_c7_3793] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l214_c2_9f76] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_cond;
     result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_return_output := result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l221_c7_3793] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l221_c7_3793_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_3793_cond;
     tmp16_MUX_uxn_opcodes_h_l221_c7_3793_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_3793_iftrue;
     tmp16_MUX_uxn_opcodes_h_l221_c7_3793_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_3793_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_3793_return_output := tmp16_MUX_uxn_opcodes_h_l221_c7_3793_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l225_c7_b145] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l221_c7_3793] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b145_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_3793_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b145_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_3793_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_b145_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_3793_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l221_c7_3793] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l221_c7_3793] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_cond;
     result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_return_output := result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l214_c2_9f76] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_cond;
     tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue;
     tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_return_output := tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l221_c7_3793] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l214_c2_9f76] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l214_c2_9f76] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_3793_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_3793_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_3793_return_output;
     REG_VAR_tmp16 := VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_9f76_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l214_c2_9f76] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_cond;
     result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_return_output := result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l214_c2_9f76] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l214_c2_9f76] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_e2b8_uxn_opcodes_h_l247_l209_DUPLICATE_d25b LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e2b8_uxn_opcodes_h_l247_l209_DUPLICATE_d25b_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_e2b8(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_9f76_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_9f76_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_9f76_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_9f76_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_9f76_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_9f76_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_9f76_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_9f76_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e2b8_uxn_opcodes_h_l247_l209_DUPLICATE_d25b_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e2b8_uxn_opcodes_h_l247_l209_DUPLICATE_d25b_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_tmp16 <= REG_VAR_tmp16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     tmp16 <= REG_COMB_tmp16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
