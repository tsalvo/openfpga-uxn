-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity sth2_0CLK_55b6500a is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sth2_0CLK_55b6500a;
architecture arch of sth2_0CLK_55b6500a is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2442_c6_d665]
signal BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2442_c2_c35c]
signal t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2442_c2_c35c]
signal t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2442_c2_c35c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2442_c2_c35c]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2442_c2_c35c]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2442_c2_c35c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2442_c2_c35c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2442_c2_c35c]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2442_c2_c35c]
signal result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2442_c2_c35c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2442_c2_c35c]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2455_c11_8016]
signal BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2455_c7_fa1f]
signal t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2455_c7_fa1f]
signal t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2455_c7_fa1f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2455_c7_fa1f]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2455_c7_fa1f]
signal result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2455_c7_fa1f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2455_c7_fa1f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2455_c7_fa1f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2458_c11_f999]
signal BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2458_c7_1494]
signal t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2458_c7_1494]
signal t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2458_c7_1494]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2458_c7_1494]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2458_c7_1494]
signal result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2458_c7_1494]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2458_c7_1494]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2458_c7_1494]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2460_c30_afd8]
signal sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2462_c11_8944]
signal BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2462_c7_a159]
signal t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2462_c7_a159]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2462_c7_a159]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2462_c7_a159]
signal result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2462_c7_a159]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2462_c7_a159]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2462_c7_a159]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2470_c11_4870]
signal BIN_OP_EQ_uxn_opcodes_h_l2470_c11_4870_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2470_c11_4870_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2470_c11_4870_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2470_c7_0fe5]
signal result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2470_c7_0fe5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2470_c7_0fe5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2470_c7_0fe5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_84a2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_vram_write := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_pc_updated := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665
BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_left,
BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_right,
BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c
t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_cond,
t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue,
t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse,
t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c
t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_cond,
t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue,
t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse,
t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c
result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c
result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c
result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c
result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c
result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c
result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016
BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_left,
BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_right,
BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f
t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond,
t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue,
t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse,
t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f
t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond,
t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue,
t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse,
t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f
result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f
result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f
result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999
BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_left,
BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_right,
BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2458_c7_1494
t16_low_MUX_uxn_opcodes_h_l2458_c7_1494 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_cond,
t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue,
t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse,
t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2458_c7_1494
t16_high_MUX_uxn_opcodes_h_l2458_c7_1494 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_cond,
t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue,
t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse,
t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494
result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494
result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_cond,
result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494
result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494
result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8
sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_ins,
sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_x,
sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_y,
sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944
BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_left,
BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_right,
BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2462_c7_a159
t16_low_MUX_uxn_opcodes_h_l2462_c7_a159 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_cond,
t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue,
t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse,
t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159
result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159
result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_cond,
result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159
result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159
result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2470_c11_4870
BIN_OP_EQ_uxn_opcodes_h_l2470_c11_4870 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2470_c11_4870_left,
BIN_OP_EQ_uxn_opcodes_h_l2470_c11_4870_right,
BIN_OP_EQ_uxn_opcodes_h_l2470_c11_4870_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5
result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_cond,
result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5
result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5
result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_return_output,
 t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output,
 t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_return_output,
 t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output,
 t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_return_output,
 t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_return_output,
 t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_return_output,
 sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_return_output,
 t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2470_c11_4870_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2442_c2_c35c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2447_c3_d0f1 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2442_c2_c35c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2452_c3_0f33 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2442_c2_c35c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2456_c3_363e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2465_c3_3715 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2467_c3_cb87 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2470_c11_4870_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2470_c11_4870_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2470_c11_4870_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2471_c3_e1f1 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2472_c3_383f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2442_l2455_l2470_l2458_DUPLICATE_7270_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2462_l2455_l2470_l2458_DUPLICATE_30d3_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2462_l2455_l2458_DUPLICATE_dc9b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2455_l2470_DUPLICATE_9c5e_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2462_l2455_l2458_DUPLICATE_9ca0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2470_l2458_DUPLICATE_7e58_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2477_l2438_DUPLICATE_69df_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_iftrue := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_right := to_unsigned(3, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2447_c3_d0f1 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2447_c3_d0f1;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2470_c11_4870_right := to_unsigned(4, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_y := resize(to_signed(-2, 3), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2452_c3_0f33 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2452_c3_0f33;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2465_c3_3715 := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2465_c3_3715;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2472_c3_383f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2472_c3_383f;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2456_c3_363e := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2456_c3_363e;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2467_c3_cb87 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2467_c3_cb87;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_right := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2471_c3_e1f1 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2471_c3_e1f1;
     VAR_sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_right := to_unsigned(2, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2470_c11_4870_left := VAR_phase;
     VAR_t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue := VAR_previous_stack_read;
     VAR_t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse := t16_high;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse := t16_low;
     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2442_l2455_l2470_l2458_DUPLICATE_7270 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2442_l2455_l2470_l2458_DUPLICATE_7270_return_output := result.u8_value;

     -- sp_relative_shift[uxn_opcodes_h_l2460_c30_afd8] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_ins;
     sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_x;
     sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_return_output := sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2442_c2_c35c] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2442_c2_c35c_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2462_l2455_l2470_l2458_DUPLICATE_30d3 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2462_l2455_l2470_l2458_DUPLICATE_30d3_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2462_l2455_l2458_DUPLICATE_9ca0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2462_l2455_l2458_DUPLICATE_9ca0_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2462_c11_8944] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_left;
     BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_return_output := BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2442_c2_c35c] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2442_c2_c35c_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2470_l2458_DUPLICATE_7e58 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2470_l2458_DUPLICATE_7e58_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2455_c11_8016] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_left;
     BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_return_output := BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2442_c6_d665] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_left;
     BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_return_output := BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2455_l2470_DUPLICATE_9c5e LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2455_l2470_DUPLICATE_9c5e_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2470_c11_4870] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2470_c11_4870_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2470_c11_4870_left;
     BIN_OP_EQ_uxn_opcodes_h_l2470_c11_4870_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2470_c11_4870_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2470_c11_4870_return_output := BIN_OP_EQ_uxn_opcodes_h_l2470_c11_4870_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2442_c2_c35c] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2442_c2_c35c_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2458_c11_f999] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_left;
     BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_return_output := BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2462_l2455_l2458_DUPLICATE_dc9b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2462_l2455_l2458_DUPLICATE_dc9b_return_output := result.is_stack_index_flipped;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2442_c6_d665_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2455_c11_8016_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2458_c11_f999_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2462_c11_8944_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2470_c11_4870_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2470_c11_4870_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2470_c11_4870_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2470_c11_4870_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2455_l2470_DUPLICATE_9c5e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2455_l2470_DUPLICATE_9c5e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2462_l2455_l2470_l2458_DUPLICATE_30d3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2462_l2455_l2470_l2458_DUPLICATE_30d3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2462_l2455_l2470_l2458_DUPLICATE_30d3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2462_l2455_l2470_l2458_DUPLICATE_30d3_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2462_l2455_l2458_DUPLICATE_dc9b_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2462_l2455_l2458_DUPLICATE_dc9b_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2462_l2455_l2458_DUPLICATE_dc9b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2462_l2455_l2458_DUPLICATE_9ca0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2462_l2455_l2458_DUPLICATE_9ca0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2462_l2455_l2458_DUPLICATE_9ca0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2470_l2458_DUPLICATE_7e58_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2470_l2458_DUPLICATE_7e58_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2442_l2455_l2470_l2458_DUPLICATE_7270_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2442_l2455_l2470_l2458_DUPLICATE_7270_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2442_l2455_l2470_l2458_DUPLICATE_7270_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2442_l2455_l2470_l2458_DUPLICATE_7270_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2442_c2_c35c_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2442_c2_c35c_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2442_c2_c35c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2460_c30_afd8_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2470_c7_0fe5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output := result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2442_c2_c35c] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2442_c2_c35c] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2462_c7_a159] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2470_c7_0fe5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2462_c7_a159] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2470_c7_0fe5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2470_c7_0fe5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2442_c2_c35c] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2462_c7_a159] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_cond;
     t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_return_output := t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2458_c7_1494] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_cond;
     t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_return_output := t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2462_c7_a159_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2462_c7_a159_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2470_c7_0fe5_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2458_c7_1494_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2462_c7_a159_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2462_c7_a159] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2462_c7_a159] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2462_c7_a159] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_return_output := result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2458_c7_1494] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_cond;
     t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_return_output := t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2458_c7_1494] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2458_c7_1494] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2462_c7_a159] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2455_c7_fa1f] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond;
     t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output := t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2462_c7_a159_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2458_c7_1494_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2458_c7_1494_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2462_c7_a159_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2462_c7_a159_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2462_c7_a159_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2458_c7_1494_return_output;
     -- t16_low_MUX[uxn_opcodes_h_l2455_c7_fa1f] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond;
     t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output := t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2458_c7_1494] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_return_output := result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2442_c2_c35c] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_cond;
     t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output := t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2455_c7_fa1f] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2458_c7_1494] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2455_c7_fa1f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2458_c7_1494] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2458_c7_1494] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2458_c7_1494_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2458_c7_1494_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2458_c7_1494_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2458_c7_1494_return_output;
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2455_c7_fa1f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2442_c2_c35c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2455_c7_fa1f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2455_c7_fa1f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2442_c2_c35c] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2455_c7_fa1f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2442_c2_c35c] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_cond;
     t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output := t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2455_c7_fa1f_return_output;
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2442_c2_c35c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2442_c2_c35c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2442_c2_c35c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2442_c2_c35c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2477_l2438_DUPLICATE_69df LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2477_l2438_DUPLICATE_69df_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_84a2(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2442_c2_c35c_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2477_l2438_DUPLICATE_69df_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2477_l2438_DUPLICATE_69df_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
