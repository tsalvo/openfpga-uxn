-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 46
entity jsr_0CLK_fedec265 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jsr_0CLK_fedec265;
architecture arch of jsr_0CLK_fedec265 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l732_c6_546c]
signal BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l732_c2_abf2]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l732_c2_abf2]
signal result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l732_c2_abf2]
signal result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l732_c2_abf2]
signal result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l732_c2_abf2]
signal result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l732_c2_abf2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l732_c2_abf2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l732_c2_abf2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_return_output : unsigned(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l732_c2_abf2]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l732_c2_abf2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l732_c2_abf2]
signal t8_MUX_uxn_opcodes_h_l732_c2_abf2_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l732_c2_abf2_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l745_c11_f793]
signal BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l745_c7_c257]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l745_c7_c257]
signal result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l745_c7_c257]
signal result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l745_c7_c257]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l745_c7_c257]
signal result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l745_c7_c257]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_return_output : unsigned(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l745_c7_c257]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l745_c7_c257]
signal result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l745_c7_c257]
signal t8_MUX_uxn_opcodes_h_l745_c7_c257_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l745_c7_c257_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l745_c7_c257_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l745_c7_c257_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l747_c30_3a46]
signal sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l749_c11_2429]
signal BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l749_c7_bd46]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l749_c7_bd46]
signal result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l749_c7_bd46]
signal result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l749_c7_bd46]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l749_c7_bd46]
signal result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l749_c7_bd46]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_return_output : unsigned(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l749_c7_bd46]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l749_c7_bd46]
signal result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l749_c7_bd46]
signal t8_MUX_uxn_opcodes_h_l749_c7_bd46_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l749_c7_bd46_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l757_c11_74b9]
signal BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l757_c7_a0e4]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l757_c7_a0e4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l757_c7_a0e4]
signal result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l757_c7_a0e4]
signal result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l757_c7_a0e4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l757_c7_a0e4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output : unsigned(0 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l760_c31_d33c]
signal CONST_SR_8_uxn_opcodes_h_l760_c31_d33c_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l760_c31_d33c_return_output : unsigned(15 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l762_c22_cbbd]
signal BIN_OP_PLUS_uxn_opcodes_h_l762_c22_cbbd_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l762_c22_cbbd_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l762_c22_cbbd_return_output : signed(17 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_500b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_pc_updated := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.u16_value := ref_toks_4;
      base.is_ram_write := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_stack_write := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_stack_index_flipped := ref_toks_9;
      base.is_opc_done := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c
BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_left,
BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_right,
BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2
result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2
result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2
result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_cond,
result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2
result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_cond,
result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2
result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2
result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2
result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2
result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_return_output);

-- t8_MUX_uxn_opcodes_h_l732_c2_abf2
t8_MUX_uxn_opcodes_h_l732_c2_abf2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l732_c2_abf2_cond,
t8_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue,
t8_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse,
t8_MUX_uxn_opcodes_h_l732_c2_abf2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793
BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_left,
BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_right,
BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257
result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257
result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_cond,
result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257
result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_cond,
result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257
result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257
result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257
result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_return_output);

-- t8_MUX_uxn_opcodes_h_l745_c7_c257
t8_MUX_uxn_opcodes_h_l745_c7_c257 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l745_c7_c257_cond,
t8_MUX_uxn_opcodes_h_l745_c7_c257_iftrue,
t8_MUX_uxn_opcodes_h_l745_c7_c257_iffalse,
t8_MUX_uxn_opcodes_h_l745_c7_c257_return_output);

-- sp_relative_shift_uxn_opcodes_h_l747_c30_3a46
sp_relative_shift_uxn_opcodes_h_l747_c30_3a46 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_ins,
sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_x,
sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_y,
sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429
BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_left,
BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_right,
BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46
result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46
result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_cond,
result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46
result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_cond,
result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46
result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46
result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46
result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_return_output);

-- t8_MUX_uxn_opcodes_h_l749_c7_bd46
t8_MUX_uxn_opcodes_h_l749_c7_bd46 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l749_c7_bd46_cond,
t8_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue,
t8_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse,
t8_MUX_uxn_opcodes_h_l749_c7_bd46_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9
BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9_left,
BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9_right,
BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4
result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4
result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4
result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_cond,
result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4
result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_cond,
result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4
result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output);

-- CONST_SR_8_uxn_opcodes_h_l760_c31_d33c
CONST_SR_8_uxn_opcodes_h_l760_c31_d33c : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l760_c31_d33c_x,
CONST_SR_8_uxn_opcodes_h_l760_c31_d33c_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l762_c22_cbbd
BIN_OP_PLUS_uxn_opcodes_h_l762_c22_cbbd : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l762_c22_cbbd_left,
BIN_OP_PLUS_uxn_opcodes_h_l762_c22_cbbd_right,
BIN_OP_PLUS_uxn_opcodes_h_l762_c22_cbbd_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_return_output,
 t8_MUX_uxn_opcodes_h_l732_c2_abf2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_return_output,
 t8_MUX_uxn_opcodes_h_l745_c7_c257_return_output,
 sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_return_output,
 t8_MUX_uxn_opcodes_h_l749_c7_bd46_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output,
 CONST_SR_8_uxn_opcodes_h_l760_c31_d33c_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l762_c22_cbbd_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l732_c2_abf2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l732_c2_abf2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l737_c3_c960 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l742_c3_4767 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l745_c7_c257_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l732_c2_abf2_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l732_c2_abf2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l746_c3_08b8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l745_c7_c257_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l745_c7_c257_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l749_c7_bd46_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l745_c7_c257_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l752_c3_253e : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l754_c3_1420 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l749_c7_bd46_cond : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l755_c21_2884_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l758_c3_47eb : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l757_c7_a0e4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l762_c3_d039 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l759_c3_54a4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l757_c7_a0e4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l760_c31_d33c_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l760_c31_d33c_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l760_c21_c53b_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l762_c22_cbbd_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l762_c27_07aa_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l762_c22_cbbd_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l762_c22_cbbd_return_output : signed(17 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l732_l757_l745_DUPLICATE_4fef_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l732_l757_l749_l745_DUPLICATE_dfab_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l757_l749_l745_DUPLICATE_97ce_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l749_l745_DUPLICATE_822b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l749_l745_DUPLICATE_ad63_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l757_l749_l745_DUPLICATE_10ad_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_500b_uxn_opcodes_h_l766_l728_DUPLICATE_d229_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l754_c3_1420 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l754_c3_1420;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l742_c3_4767 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l742_c3_4767;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l752_c3_253e := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l752_c3_253e;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_right := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l737_c3_c960 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l737_c3_c960;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l759_c3_54a4 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l759_c3_54a4;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9_right := to_unsigned(3, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l746_c3_08b8 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l746_c3_08b8;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l758_c3_47eb := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l758_c3_47eb;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_ins := VAR_ins;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l762_c22_cbbd_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_CONST_SR_8_uxn_opcodes_h_l760_c31_d33c_x := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l745_c7_c257_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l757_c11_74b9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9_left;
     BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9_return_output := BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l732_c2_abf2] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l732_c2_abf2_return_output := result.is_vram_write;

     -- result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d[uxn_opcodes_h_l757_c7_a0e4] LATENCY=0
     VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l757_c7_a0e4_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l757_l749_l745_DUPLICATE_10ad LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l757_l749_l745_DUPLICATE_10ad_return_output := result.is_opc_done;

     -- sp_relative_shift[uxn_opcodes_h_l747_c30_3a46] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_ins;
     sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_x <= VAR_sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_x;
     sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_y <= VAR_sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_return_output := sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l732_c2_abf2] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l732_c2_abf2_return_output := result.is_ram_write;

     -- CAST_TO_int8_t[uxn_opcodes_h_l762_c27_07aa] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l762_c27_07aa_return_output := CAST_TO_int8_t_uint8_t(
     t8);

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l749_l745_DUPLICATE_ad63 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l749_l745_DUPLICATE_ad63_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l732_l757_l749_l745_DUPLICATE_dfab LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l732_l757_l749_l745_DUPLICATE_dfab_return_output := result.u16_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l732_c6_546c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_left;
     BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_return_output := BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l732_l757_l745_DUPLICATE_4fef LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l732_l757_l745_DUPLICATE_4fef_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l745_c11_f793] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_left;
     BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_return_output := BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_return_output;

     -- CONST_SR_8[uxn_opcodes_h_l760_c31_d33c] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l760_c31_d33c_x <= VAR_CONST_SR_8_uxn_opcodes_h_l760_c31_d33c_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l760_c31_d33c_return_output := CONST_SR_8_uxn_opcodes_h_l760_c31_d33c_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l757_l749_l745_DUPLICATE_97ce LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l757_l749_l745_DUPLICATE_97ce_return_output := result.is_pc_updated;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l757_c7_a0e4] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l757_c7_a0e4_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l749_c11_2429] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_left;
     BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_return_output := BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l749_l745_DUPLICATE_822b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l749_l745_DUPLICATE_822b_return_output := result.is_stack_write;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l755_c21_2884] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l755_c21_2884_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_pc);

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l732_c2_abf2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c6_546c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l745_c7_c257_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l745_c11_f793_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l749_c7_bd46_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_2429_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l757_c11_74b9_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l762_c22_cbbd_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l762_c27_07aa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l755_c21_2884_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l732_l757_l749_l745_DUPLICATE_dfab_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l732_l757_l749_l745_DUPLICATE_dfab_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l732_l757_l749_l745_DUPLICATE_dfab_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l732_l757_l749_l745_DUPLICATE_dfab_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l757_l749_l745_DUPLICATE_10ad_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l757_l749_l745_DUPLICATE_10ad_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l757_l749_l745_DUPLICATE_10ad_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l757_l749_l745_DUPLICATE_97ce_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l757_l749_l745_DUPLICATE_97ce_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l757_l749_l745_DUPLICATE_97ce_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l749_l745_DUPLICATE_ad63_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l749_l745_DUPLICATE_ad63_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l749_l745_DUPLICATE_822b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l749_l745_DUPLICATE_822b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l732_l757_l745_DUPLICATE_4fef_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l732_l757_l745_DUPLICATE_4fef_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l732_l757_l745_DUPLICATE_4fef_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l732_c2_abf2_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l732_c2_abf2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse := VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l757_c7_a0e4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l757_c7_a0e4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l747_c30_3a46_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l757_c7_a0e4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l732_c2_abf2] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l762_c22_cbbd] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l762_c22_cbbd_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l762_c22_cbbd_left;
     BIN_OP_PLUS_uxn_opcodes_h_l762_c22_cbbd_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l762_c22_cbbd_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l762_c22_cbbd_return_output := BIN_OP_PLUS_uxn_opcodes_h_l762_c22_cbbd_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l749_c7_bd46] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l760_c21_c53b] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l760_c21_c53b_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l760_c31_d33c_return_output);

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l757_c7_a0e4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l757_c7_a0e4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l732_c2_abf2] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l749_c7_bd46] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l757_c7_a0e4] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output;

     -- t8_MUX[uxn_opcodes_h_l749_c7_bd46] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l749_c7_bd46_cond <= VAR_t8_MUX_uxn_opcodes_h_l749_c7_bd46_cond;
     t8_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue;
     t8_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l749_c7_bd46_return_output := t8_MUX_uxn_opcodes_h_l749_c7_bd46_return_output;

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l762_c3_d039 := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l762_c22_cbbd_return_output)),16);
     VAR_result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l760_c21_c53b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_bd46_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_bd46_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l745_c7_c257_iffalse := VAR_t8_MUX_uxn_opcodes_h_l749_c7_bd46_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue := VAR_result_u16_value_uxn_opcodes_h_l762_c3_d039;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l749_c7_bd46] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l745_c7_c257] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l745_c7_c257] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l749_c7_bd46] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l749_c7_bd46] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_return_output;

     -- t8_MUX[uxn_opcodes_h_l745_c7_c257] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l745_c7_c257_cond <= VAR_t8_MUX_uxn_opcodes_h_l745_c7_c257_cond;
     t8_MUX_uxn_opcodes_h_l745_c7_c257_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l745_c7_c257_iftrue;
     t8_MUX_uxn_opcodes_h_l745_c7_c257_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l745_c7_c257_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l745_c7_c257_return_output := t8_MUX_uxn_opcodes_h_l745_c7_c257_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l757_c7_a0e4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output := result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l749_c7_bd46] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l757_c7_a0e4] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_cond;
     result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output := result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_bd46_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_bd46_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l745_c7_c257_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l745_c7_c257_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_bd46_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_bd46_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l757_c7_a0e4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse := VAR_t8_MUX_uxn_opcodes_h_l745_c7_c257_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l745_c7_c257] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_return_output;

     -- t8_MUX[uxn_opcodes_h_l732_c2_abf2] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l732_c2_abf2_cond <= VAR_t8_MUX_uxn_opcodes_h_l732_c2_abf2_cond;
     t8_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue;
     t8_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l732_c2_abf2_return_output := t8_MUX_uxn_opcodes_h_l732_c2_abf2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l732_c2_abf2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l732_c2_abf2] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l749_c7_bd46] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_cond;
     result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_return_output := result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l745_c7_c257] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l745_c7_c257] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l745_c7_c257] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l749_c7_bd46] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_cond;
     result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_return_output := result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l745_c7_c257_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l745_c7_c257_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l745_c7_c257_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l745_c7_c257_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c7_bd46_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l749_c7_bd46_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l732_c2_abf2_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l745_c7_c257] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_cond;
     result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_return_output := result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l732_c2_abf2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l745_c7_c257] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_cond;
     result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_return_output := result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l732_c2_abf2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l732_c2_abf2] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l732_c2_abf2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_return_output;

     -- Submodule level 5
     VAR_result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l745_c7_c257_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l745_c7_c257_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l732_c2_abf2] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_cond;
     result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_return_output := result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l732_c2_abf2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_return_output := result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_500b_uxn_opcodes_h_l766_l728_DUPLICATE_d229 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_500b_uxn_opcodes_h_l766_l728_DUPLICATE_d229_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_500b(
     result,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l732_c2_abf2_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l732_c2_abf2_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l732_c2_abf2_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l732_c2_abf2_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l732_c2_abf2_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l732_c2_abf2_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l732_c2_abf2_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c2_abf2_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c2_abf2_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l732_c2_abf2_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_500b_uxn_opcodes_h_l766_l728_DUPLICATE_d229_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_500b_uxn_opcodes_h_l766_l728_DUPLICATE_d229_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
