-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 29
entity sth_0CLK_a9f1e08f is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sth_0CLK_a9f1e08f;
architecture arch of sth_0CLK_a9f1e08f is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2409_c6_e540]
signal BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2409_c2_cab1]
signal t8_MUX_uxn_opcodes_h_l2409_c2_cab1_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2409_c2_cab1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2409_c2_cab1]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2409_c2_cab1]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2409_c2_cab1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2409_c2_cab1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2409_c2_cab1]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2409_c2_cab1]
signal result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2409_c2_cab1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2409_c2_cab1]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2422_c11_dd7f]
signal BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2422_c7_f4db]
signal t8_MUX_uxn_opcodes_h_l2422_c7_f4db_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2422_c7_f4db]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2422_c7_f4db]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2422_c7_f4db]
signal result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2422_c7_f4db]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2422_c7_f4db]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2422_c7_f4db]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2423_c30_a5f7]
signal sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2425_c11_7a9b]
signal BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2425_c7_e433]
signal t8_MUX_uxn_opcodes_h_l2425_c7_e433_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2425_c7_e433_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2425_c7_e433]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2425_c7_e433]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2425_c7_e433]
signal result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2425_c7_e433]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2425_c7_e433]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2425_c7_e433]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_84a2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_vram_write := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_pc_updated := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540
BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_left,
BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_right,
BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_return_output);

-- t8_MUX_uxn_opcodes_h_l2409_c2_cab1
t8_MUX_uxn_opcodes_h_l2409_c2_cab1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2409_c2_cab1_cond,
t8_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue,
t8_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse,
t8_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1
result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1
result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1
result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1
result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1
result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1
result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_cond,
result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1
result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f
BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_left,
BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_right,
BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_return_output);

-- t8_MUX_uxn_opcodes_h_l2422_c7_f4db
t8_MUX_uxn_opcodes_h_l2422_c7_f4db : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2422_c7_f4db_cond,
t8_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue,
t8_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse,
t8_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db
result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db
result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_cond,
result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db
result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db
result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7
sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_ins,
sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_x,
sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_y,
sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b
BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_left,
BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_right,
BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_return_output);

-- t8_MUX_uxn_opcodes_h_l2425_c7_e433
t8_MUX_uxn_opcodes_h_l2425_c7_e433 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2425_c7_e433_cond,
t8_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue,
t8_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse,
t8_MUX_uxn_opcodes_h_l2425_c7_e433_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433
result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_cond,
result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433
result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_return_output,
 t8_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_return_output,
 t8_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output,
 sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_return_output,
 t8_MUX_uxn_opcodes_h_l2425_c7_e433_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2409_c2_cab1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2409_c2_cab1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2414_c3_d600 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2409_c2_cab1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2419_c3_fa8a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2409_c2_cab1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2425_c7_e433_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2422_c7_f4db_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2425_c7_e433_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2428_c3_0716 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2425_c7_e433_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2430_c3_1f2c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2409_l2422_l2425_DUPLICATE_26e9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2422_l2425_DUPLICATE_504d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2422_l2425_DUPLICATE_bf38_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2422_l2425_DUPLICATE_0441_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2422_l2425_DUPLICATE_7cc0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2435_l2405_DUPLICATE_7cb8_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2428_c3_0716 := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2428_c3_0716;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2419_c3_fa8a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2419_c3_fa8a;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2414_c3_d600 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2414_c3_d600;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2430_c3_1f2c := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2430_c3_1f2c;
     VAR_sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_right := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2422_c11_dd7f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2423_c30_a5f7] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_ins;
     sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_x;
     sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_return_output := sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_return_output;

     -- result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d[uxn_opcodes_h_l2425_c7_e433] LATENCY=0
     VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2425_c7_e433_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2422_l2425_DUPLICATE_504d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2422_l2425_DUPLICATE_504d_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2409_c6_e540] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_left;
     BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_return_output := BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2409_c2_cab1] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2409_c2_cab1_return_output := result.is_vram_write;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2409_c2_cab1] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2409_c2_cab1_return_output := result.is_ram_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2409_c2_cab1] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2409_c2_cab1_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l2425_c11_7a9b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_left;
     BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_return_output := BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2422_l2425_DUPLICATE_bf38 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2422_l2425_DUPLICATE_bf38_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2422_l2425_DUPLICATE_7cc0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2422_l2425_DUPLICATE_7cc0_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2422_l2425_DUPLICATE_0441 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2422_l2425_DUPLICATE_0441_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2409_l2422_l2425_DUPLICATE_26e9 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2409_l2422_l2425_DUPLICATE_26e9_return_output := result.u8_value;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2409_c2_cab1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2409_c6_e540_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2422_c7_f4db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_dd7f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2425_c7_e433_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_7a9b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2422_l2425_DUPLICATE_504d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2422_l2425_DUPLICATE_504d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2422_l2425_DUPLICATE_bf38_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2422_l2425_DUPLICATE_bf38_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2422_l2425_DUPLICATE_7cc0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2422_l2425_DUPLICATE_7cc0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2422_l2425_DUPLICATE_0441_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2422_l2425_DUPLICATE_0441_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2409_l2422_l2425_DUPLICATE_26e9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2409_l2422_l2425_DUPLICATE_26e9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2409_l2422_l2425_DUPLICATE_26e9_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2409_c2_cab1_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2409_c2_cab1_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2409_c2_cab1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse := VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2425_c7_e433_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2423_c30_a5f7_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2425_c7_e433] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_return_output;

     -- t8_MUX[uxn_opcodes_h_l2425_c7_e433] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2425_c7_e433_cond <= VAR_t8_MUX_uxn_opcodes_h_l2425_c7_e433_cond;
     t8_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue;
     t8_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2425_c7_e433_return_output := t8_MUX_uxn_opcodes_h_l2425_c7_e433_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2425_c7_e433] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2409_c2_cab1] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2425_c7_e433] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2425_c7_e433] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2425_c7_e433] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2425_c7_e433] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_return_output := result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2409_c2_cab1] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2409_c2_cab1] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_e433_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2425_c7_e433_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_e433_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_e433_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_e433_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_e433_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2425_c7_e433_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2422_c7_f4db] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2422_c7_f4db] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2422_c7_f4db] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output;

     -- t8_MUX[uxn_opcodes_h_l2422_c7_f4db] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2422_c7_f4db_cond <= VAR_t8_MUX_uxn_opcodes_h_l2422_c7_f4db_cond;
     t8_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue;
     t8_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output := t8_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2422_c7_f4db] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output := result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2422_c7_f4db] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2422_c7_f4db] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2422_c7_f4db_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2409_c2_cab1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2409_c2_cab1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output := result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2409_c2_cab1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2409_c2_cab1] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output;

     -- t8_MUX[uxn_opcodes_h_l2409_c2_cab1] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2409_c2_cab1_cond <= VAR_t8_MUX_uxn_opcodes_h_l2409_c2_cab1_cond;
     t8_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue;
     t8_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output := t8_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2409_c2_cab1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2409_c2_cab1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output;

     -- Submodule level 4
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2435_l2405_DUPLICATE_7cb8 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2435_l2405_DUPLICATE_7cb8_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_84a2(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2409_c2_cab1_return_output);

     -- Submodule level 5
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2435_l2405_DUPLICATE_7cb8_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2435_l2405_DUPLICATE_7cb8_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
