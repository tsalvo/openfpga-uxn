-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 47
entity dup_0CLK_a148083c is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dup_0CLK_a148083c;
architecture arch of dup_0CLK_a148083c is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l3153_c6_ddae]
signal BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l3153_c1_e760]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l3153_c2_5808]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_return_output : unsigned(0 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l3153_c2_5808]
signal result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l3153_c2_5808]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l3153_c2_5808]
signal result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3153_c2_5808]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l3153_c2_5808]
signal result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l3153_c2_5808]
signal result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l3153_c2_5808]
signal t8_MUX_uxn_opcodes_h_l3153_c2_5808_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l3153_c2_5808_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l3154_c3_7477[uxn_opcodes_h_l3154_c3_7477]
signal printf_uxn_opcodes_h_l3154_c3_7477_uxn_opcodes_h_l3154_c3_7477_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l3159_c11_6546]
signal BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l3159_c7_9247]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_return_output : unsigned(0 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l3159_c7_9247]
signal result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l3159_c7_9247]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l3159_c7_9247]
signal result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3159_c7_9247]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l3159_c7_9247]
signal result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l3159_c7_9247]
signal result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l3159_c7_9247]
signal t8_MUX_uxn_opcodes_h_l3159_c7_9247_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l3159_c7_9247_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l3162_c11_16e2]
signal BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l3162_c7_a6da]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output : unsigned(0 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l3162_c7_a6da]
signal result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l3162_c7_a6da]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l3162_c7_a6da]
signal result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3162_c7_a6da]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l3162_c7_a6da]
signal result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l3162_c7_a6da]
signal result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l3162_c7_a6da]
signal t8_MUX_uxn_opcodes_h_l3162_c7_a6da_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output : unsigned(7 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l3166_c32_96aa]
signal BIN_OP_AND_uxn_opcodes_h_l3166_c32_96aa_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l3166_c32_96aa_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l3166_c32_96aa_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l3166_c32_6088]
signal BIN_OP_GT_uxn_opcodes_h_l3166_c32_6088_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l3166_c32_6088_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l3166_c32_6088_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l3166_c32_6c09]
signal MUX_uxn_opcodes_h_l3166_c32_6c09_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l3166_c32_6c09_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l3166_c32_6c09_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l3166_c32_6c09_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l3168_c11_8fd0]
signal BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l3168_c7_db6f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l3168_c7_db6f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l3168_c7_db6f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3168_c7_db6f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l3168_c7_db6f]
signal result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l3174_c11_5a4f]
signal BIN_OP_EQ_uxn_opcodes_h_l3174_c11_5a4f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3174_c11_5a4f_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3174_c11_5a4f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l3174_c7_5393]
signal result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l3174_c7_5393]
signal result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3174_c7_5393]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l3174_c7_5393]
signal result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l3178_c11_9237]
signal BIN_OP_EQ_uxn_opcodes_h_l3178_c11_9237_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3178_c11_9237_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l3178_c11_9237_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l3178_c7_0262]
signal result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l3178_c7_0262]
signal result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_1ade( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_sp_shift := ref_toks_1;
      base.is_stack_read := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_opc_done := ref_toks_6;
      base.stack_value := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae
BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_left,
BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_right,
BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808
result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808
result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808
result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808
result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808
result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808
result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_cond,
result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_return_output);

-- t8_MUX_uxn_opcodes_h_l3153_c2_5808
t8_MUX_uxn_opcodes_h_l3153_c2_5808 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l3153_c2_5808_cond,
t8_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue,
t8_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse,
t8_MUX_uxn_opcodes_h_l3153_c2_5808_return_output);

-- printf_uxn_opcodes_h_l3154_c3_7477_uxn_opcodes_h_l3154_c3_7477
printf_uxn_opcodes_h_l3154_c3_7477_uxn_opcodes_h_l3154_c3_7477 : entity work.printf_uxn_opcodes_h_l3154_c3_7477_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l3154_c3_7477_uxn_opcodes_h_l3154_c3_7477_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546
BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_left,
BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_right,
BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247
result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247
result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247
result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247
result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247
result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247
result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_cond,
result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_return_output);

-- t8_MUX_uxn_opcodes_h_l3159_c7_9247
t8_MUX_uxn_opcodes_h_l3159_c7_9247 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l3159_c7_9247_cond,
t8_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue,
t8_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse,
t8_MUX_uxn_opcodes_h_l3159_c7_9247_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2
BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_left,
BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_right,
BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da
result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da
result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da
result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da
result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da
result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da
result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_cond,
result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output);

-- t8_MUX_uxn_opcodes_h_l3162_c7_a6da
t8_MUX_uxn_opcodes_h_l3162_c7_a6da : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l3162_c7_a6da_cond,
t8_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue,
t8_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse,
t8_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l3166_c32_96aa
BIN_OP_AND_uxn_opcodes_h_l3166_c32_96aa : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l3166_c32_96aa_left,
BIN_OP_AND_uxn_opcodes_h_l3166_c32_96aa_right,
BIN_OP_AND_uxn_opcodes_h_l3166_c32_96aa_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l3166_c32_6088
BIN_OP_GT_uxn_opcodes_h_l3166_c32_6088 : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l3166_c32_6088_left,
BIN_OP_GT_uxn_opcodes_h_l3166_c32_6088_right,
BIN_OP_GT_uxn_opcodes_h_l3166_c32_6088_return_output);

-- MUX_uxn_opcodes_h_l3166_c32_6c09
MUX_uxn_opcodes_h_l3166_c32_6c09 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l3166_c32_6c09_cond,
MUX_uxn_opcodes_h_l3166_c32_6c09_iftrue,
MUX_uxn_opcodes_h_l3166_c32_6c09_iffalse,
MUX_uxn_opcodes_h_l3166_c32_6c09_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0
BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0_left,
BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0_right,
BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f
result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f
result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f
result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f
result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_cond,
result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l3174_c11_5a4f
BIN_OP_EQ_uxn_opcodes_h_l3174_c11_5a4f : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l3174_c11_5a4f_left,
BIN_OP_EQ_uxn_opcodes_h_l3174_c11_5a4f_right,
BIN_OP_EQ_uxn_opcodes_h_l3174_c11_5a4f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393
result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393
result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393
result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_cond,
result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l3178_c11_9237
BIN_OP_EQ_uxn_opcodes_h_l3178_c11_9237 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l3178_c11_9237_left,
BIN_OP_EQ_uxn_opcodes_h_l3178_c11_9237_right,
BIN_OP_EQ_uxn_opcodes_h_l3178_c11_9237_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262
result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262
result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_return_output,
 t8_MUX_uxn_opcodes_h_l3153_c2_5808_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_return_output,
 t8_MUX_uxn_opcodes_h_l3159_c7_9247_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output,
 t8_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output,
 BIN_OP_AND_uxn_opcodes_h_l3166_c32_96aa_return_output,
 BIN_OP_GT_uxn_opcodes_h_l3166_c32_6088_return_output,
 MUX_uxn_opcodes_h_l3166_c32_6c09_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l3174_c11_5a4f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l3178_c11_9237_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3156_c3_6088 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3159_c7_9247_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3153_c2_5808_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3153_c2_5808_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l3154_c3_7477_uxn_opcodes_h_l3154_c3_7477_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3160_c3_6dc0 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3159_c7_9247_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l3162_c7_a6da_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l3166_c32_6c09_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l3166_c32_6c09_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l3166_c32_6c09_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l3166_c32_96aa_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l3166_c32_96aa_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l3166_c32_96aa_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l3166_c32_6088_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l3166_c32_6088_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l3166_c32_6088_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l3166_c32_6c09_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3171_c3_53b3 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3174_c11_5a4f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3174_c11_5a4f_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3174_c11_5a4f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3175_c3_1dda : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3178_c11_9237_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3178_c11_9237_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l3178_c11_9237_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l3168_l3159_l3153_DUPLICATE_51ae_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l3159_l3162_l3153_DUPLICATE_fe05_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3159_l3153_l3178_l3174_l3162_DUPLICATE_1f1f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3159_l3174_l3162_l3153_DUPLICATE_0995_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l3159_l3162_DUPLICATE_bc3e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3159_l3178_l3174_l3168_l3162_DUPLICATE_6e61_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l3174_l3162_DUPLICATE_6e19_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1ade_uxn_opcodes_h_l3183_l3149_DUPLICATE_490b_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_GT_uxn_opcodes_h_l3166_c32_6088_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_right := to_unsigned(2, 2);
     VAR_MUX_uxn_opcodes_h_l3166_c32_6c09_iffalse := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3171_c3_53b3 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3171_c3_53b3;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_iftrue := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3156_c3_6088 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3156_c3_6088;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3174_c11_5a4f_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3178_c11_9237_right := to_unsigned(5, 3);
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3175_c3_1dda := resize(to_unsigned(2, 2), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3175_c3_1dda;
     VAR_MUX_uxn_opcodes_h_l3166_c32_6c09_iftrue := signed(std_logic_vector(resize(to_unsigned(2, 2), 8)));
     VAR_BIN_OP_AND_uxn_opcodes_h_l3166_c32_96aa_right := to_unsigned(128, 8);
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3160_c3_6dc0 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l3160_c3_6dc0;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_AND_uxn_opcodes_h_l3166_c32_96aa_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3174_c11_5a4f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3178_c11_9237_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue := VAR_previous_stack_read;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue := t8;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3159_l3153_l3178_l3174_l3162_DUPLICATE_1f1f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3159_l3153_l3178_l3174_l3162_DUPLICATE_1f1f_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l3153_c6_ddae] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_left;
     BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_return_output := BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l3159_c11_6546] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_left;
     BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_return_output := BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3159_l3174_l3162_l3153_DUPLICATE_0995 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3159_l3174_l3162_l3153_DUPLICATE_0995_return_output := result.stack_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l3168_l3159_l3153_DUPLICATE_51ae LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l3168_l3159_l3153_DUPLICATE_51ae_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l3174_l3162_DUPLICATE_6e19 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l3174_l3162_DUPLICATE_6e19_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l3162_c11_16e2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_left;
     BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_return_output := BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l3166_c32_96aa] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l3166_c32_96aa_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l3166_c32_96aa_left;
     BIN_OP_AND_uxn_opcodes_h_l3166_c32_96aa_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l3166_c32_96aa_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l3166_c32_96aa_return_output := BIN_OP_AND_uxn_opcodes_h_l3166_c32_96aa_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l3159_l3162_DUPLICATE_bc3e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l3159_l3162_DUPLICATE_bc3e_return_output := result.is_stack_read;

     -- BIN_OP_EQ[uxn_opcodes_h_l3178_c11_9237] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l3178_c11_9237_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3178_c11_9237_left;
     BIN_OP_EQ_uxn_opcodes_h_l3178_c11_9237_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3178_c11_9237_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3178_c11_9237_return_output := BIN_OP_EQ_uxn_opcodes_h_l3178_c11_9237_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l3174_c11_5a4f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l3174_c11_5a4f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3174_c11_5a4f_left;
     BIN_OP_EQ_uxn_opcodes_h_l3174_c11_5a4f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3174_c11_5a4f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3174_c11_5a4f_return_output := BIN_OP_EQ_uxn_opcodes_h_l3174_c11_5a4f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l3168_c11_8fd0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0_left;
     BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0_return_output := BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0_return_output;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l3159_l3162_l3153_DUPLICATE_fe05 LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l3159_l3162_l3153_DUPLICATE_fe05_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3159_l3178_l3174_l3168_l3162_DUPLICATE_6e61 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3159_l3178_l3174_l3168_l3162_DUPLICATE_6e61_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l3166_c32_6088_left := VAR_BIN_OP_AND_uxn_opcodes_h_l3166_c32_96aa_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l3153_c2_5808_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3153_c6_ddae_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l3159_c7_9247_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3159_c11_6546_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l3162_c7_a6da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3162_c11_16e2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3168_c11_8fd0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3174_c11_5a4f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3174_c11_5a4f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3174_c11_5a4f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3174_c11_5a4f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3178_c11_9237_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l3178_c11_9237_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l3159_l3162_l3153_DUPLICATE_fe05_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l3159_l3162_l3153_DUPLICATE_fe05_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l3159_l3162_l3153_DUPLICATE_fe05_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3159_l3178_l3174_l3168_l3162_DUPLICATE_6e61_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3159_l3178_l3174_l3168_l3162_DUPLICATE_6e61_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3159_l3178_l3174_l3168_l3162_DUPLICATE_6e61_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3159_l3178_l3174_l3168_l3162_DUPLICATE_6e61_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l3159_l3178_l3174_l3168_l3162_DUPLICATE_6e61_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l3168_l3159_l3153_DUPLICATE_51ae_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l3168_l3159_l3153_DUPLICATE_51ae_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l3168_l3159_l3153_DUPLICATE_51ae_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l3159_l3162_DUPLICATE_bc3e_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l3159_l3162_DUPLICATE_bc3e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3159_l3153_l3178_l3174_l3162_DUPLICATE_1f1f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3159_l3153_l3178_l3174_l3162_DUPLICATE_1f1f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3159_l3153_l3178_l3174_l3162_DUPLICATE_1f1f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3159_l3153_l3178_l3174_l3162_DUPLICATE_1f1f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l3159_l3153_l3178_l3174_l3162_DUPLICATE_1f1f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l3174_l3162_DUPLICATE_6e19_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l3174_l3162_DUPLICATE_6e19_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3159_l3174_l3162_l3153_DUPLICATE_0995_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3159_l3174_l3162_l3153_DUPLICATE_0995_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3159_l3174_l3162_l3153_DUPLICATE_0995_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l3159_l3174_l3162_l3153_DUPLICATE_0995_return_output;
     -- BIN_OP_GT[uxn_opcodes_h_l3166_c32_6088] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l3166_c32_6088_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l3166_c32_6088_left;
     BIN_OP_GT_uxn_opcodes_h_l3166_c32_6088_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l3166_c32_6088_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l3166_c32_6088_return_output := BIN_OP_GT_uxn_opcodes_h_l3166_c32_6088_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l3178_c7_0262] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l3174_c7_5393] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_cond;
     result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_return_output := result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l3162_c7_a6da] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l3178_c7_0262] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_return_output;

     -- t8_MUX[uxn_opcodes_h_l3162_c7_a6da] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l3162_c7_a6da_cond <= VAR_t8_MUX_uxn_opcodes_h_l3162_c7_a6da_cond;
     t8_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue;
     t8_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output := t8_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l3168_c7_db6f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l3153_c1_e760] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3174_c7_5393] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l3166_c32_6c09_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l3166_c32_6088_return_output;
     VAR_printf_uxn_opcodes_h_l3154_c3_7477_uxn_opcodes_h_l3154_c3_7477_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l3153_c1_e760_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3178_c7_0262_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3178_c7_0262_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3174_c7_5393_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l3174_c7_5393_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse := VAR_t8_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l3162_c7_a6da] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output;

     -- printf_uxn_opcodes_h_l3154_c3_7477[uxn_opcodes_h_l3154_c3_7477] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l3154_c3_7477_uxn_opcodes_h_l3154_c3_7477_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l3154_c3_7477_uxn_opcodes_h_l3154_c3_7477_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- MUX[uxn_opcodes_h_l3166_c32_6c09] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l3166_c32_6c09_cond <= VAR_MUX_uxn_opcodes_h_l3166_c32_6c09_cond;
     MUX_uxn_opcodes_h_l3166_c32_6c09_iftrue <= VAR_MUX_uxn_opcodes_h_l3166_c32_6c09_iftrue;
     MUX_uxn_opcodes_h_l3166_c32_6c09_iffalse <= VAR_MUX_uxn_opcodes_h_l3166_c32_6c09_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l3166_c32_6c09_return_output := MUX_uxn_opcodes_h_l3166_c32_6c09_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l3174_c7_5393] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_return_output;

     -- t8_MUX[uxn_opcodes_h_l3159_c7_9247] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l3159_c7_9247_cond <= VAR_t8_MUX_uxn_opcodes_h_l3159_c7_9247_cond;
     t8_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue;
     t8_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l3159_c7_9247_return_output := t8_MUX_uxn_opcodes_h_l3159_c7_9247_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l3174_c7_5393] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l3159_c7_9247] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l3168_c7_db6f] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_cond;
     result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output := result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3168_c7_db6f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue := VAR_MUX_uxn_opcodes_h_l3166_c32_6c09_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3174_c7_5393_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3159_c7_9247_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3174_c7_5393_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse := VAR_t8_MUX_uxn_opcodes_h_l3159_c7_9247_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3162_c7_a6da] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l3162_c7_a6da] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_cond;
     result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output := result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l3168_c7_db6f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l3162_c7_a6da] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l3168_c7_db6f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output;

     -- t8_MUX[uxn_opcodes_h_l3153_c2_5808] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l3153_c2_5808_cond <= VAR_t8_MUX_uxn_opcodes_h_l3153_c2_5808_cond;
     t8_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue;
     t8_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l3153_c2_5808_return_output := t8_MUX_uxn_opcodes_h_l3153_c2_5808_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l3159_c7_9247] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l3153_c2_5808] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3159_c7_9247_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3168_c7_db6f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l3153_c2_5808_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3159_c7_9247] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l3159_c7_9247] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l3159_c7_9247] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_cond;
     result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_return_output := result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l3153_c2_5808] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l3162_c7_a6da] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l3162_c7_a6da] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3162_c7_a6da_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3159_c7_9247_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3159_c7_9247_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l3159_c7_9247_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l3159_c7_9247] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l3153_c2_5808] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_cond;
     result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_return_output := result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l3153_c2_5808] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l3159_c7_9247] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l3153_c2_5808] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3159_c7_9247_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3159_c7_9247_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l3153_c2_5808] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l3153_c2_5808] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_1ade_uxn_opcodes_h_l3183_l3149_DUPLICATE_490b LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1ade_uxn_opcodes_h_l3183_l3149_DUPLICATE_490b_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_1ade(
     result,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l3153_c2_5808_return_output,
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l3153_c2_5808_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l3153_c2_5808_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l3153_c2_5808_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l3153_c2_5808_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l3153_c2_5808_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l3153_c2_5808_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1ade_uxn_opcodes_h_l3183_l3149_DUPLICATE_490b_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1ade_uxn_opcodes_h_l3183_l3149_DUPLICATE_490b_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
