-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity neq_0CLK_85d5529e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end neq_0CLK_85d5529e;
architecture arch of neq_0CLK_85d5529e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1188_c6_a30b]
signal BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1188_c1_1dc7]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1188_c2_a4da]
signal n8_MUX_uxn_opcodes_h_l1188_c2_a4da_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1188_c2_a4da]
signal t8_MUX_uxn_opcodes_h_l1188_c2_a4da_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1188_c2_a4da]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1188_c2_a4da]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1188_c2_a4da]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1188_c2_a4da]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1188_c2_a4da]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1188_c2_a4da]
signal result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1189_c3_7acb[uxn_opcodes_h_l1189_c3_7acb]
signal printf_uxn_opcodes_h_l1189_c3_7acb_uxn_opcodes_h_l1189_c3_7acb_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1193_c11_c6fc]
signal BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1193_c7_cbcd]
signal n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1193_c7_cbcd]
signal t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1193_c7_cbcd]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1193_c7_cbcd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1193_c7_cbcd]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1193_c7_cbcd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1193_c7_cbcd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1193_c7_cbcd]
signal result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1196_c11_4891]
signal BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1196_c7_43ef]
signal n8_MUX_uxn_opcodes_h_l1196_c7_43ef_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1196_c7_43ef]
signal t8_MUX_uxn_opcodes_h_l1196_c7_43ef_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1196_c7_43ef]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1196_c7_43ef]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1196_c7_43ef]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1196_c7_43ef]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1196_c7_43ef]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1196_c7_43ef]
signal result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1199_c11_f09c]
signal BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1199_c7_28f4]
signal n8_MUX_uxn_opcodes_h_l1199_c7_28f4_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1199_c7_28f4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1199_c7_28f4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1199_c7_28f4]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1199_c7_28f4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1199_c7_28f4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1199_c7_28f4]
signal result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1202_c30_11fe]
signal sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1205_c21_4630]
signal BIN_OP_EQ_uxn_opcodes_h_l1205_c21_4630_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1205_c21_4630_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1205_c21_4630_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1205_c21_c121]
signal MUX_uxn_opcodes_h_l1205_c21_c121_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1205_c21_c121_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1205_c21_c121_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1205_c21_c121_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1207_c11_acd0]
signal BIN_OP_EQ_uxn_opcodes_h_l1207_c11_acd0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1207_c11_acd0_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1207_c11_acd0_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1207_c7_46ff]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1207_c7_46ff]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1207_c7_46ff]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_5b93( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b
BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_left,
BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_right,
BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_return_output);

-- n8_MUX_uxn_opcodes_h_l1188_c2_a4da
n8_MUX_uxn_opcodes_h_l1188_c2_a4da : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1188_c2_a4da_cond,
n8_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue,
n8_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse,
n8_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output);

-- t8_MUX_uxn_opcodes_h_l1188_c2_a4da
t8_MUX_uxn_opcodes_h_l1188_c2_a4da : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1188_c2_a4da_cond,
t8_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue,
t8_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse,
t8_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da
result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da
result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da
result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da
result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da
result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_cond,
result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output);

-- printf_uxn_opcodes_h_l1189_c3_7acb_uxn_opcodes_h_l1189_c3_7acb
printf_uxn_opcodes_h_l1189_c3_7acb_uxn_opcodes_h_l1189_c3_7acb : entity work.printf_uxn_opcodes_h_l1189_c3_7acb_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1189_c3_7acb_uxn_opcodes_h_l1189_c3_7acb_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc
BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_left,
BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_right,
BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_return_output);

-- n8_MUX_uxn_opcodes_h_l1193_c7_cbcd
n8_MUX_uxn_opcodes_h_l1193_c7_cbcd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond,
n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue,
n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse,
n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output);

-- t8_MUX_uxn_opcodes_h_l1193_c7_cbcd
t8_MUX_uxn_opcodes_h_l1193_c7_cbcd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond,
t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue,
t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse,
t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd
result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd
result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd
result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd
result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd
result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond,
result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891
BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_left,
BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_right,
BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_return_output);

-- n8_MUX_uxn_opcodes_h_l1196_c7_43ef
n8_MUX_uxn_opcodes_h_l1196_c7_43ef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1196_c7_43ef_cond,
n8_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue,
n8_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse,
n8_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output);

-- t8_MUX_uxn_opcodes_h_l1196_c7_43ef
t8_MUX_uxn_opcodes_h_l1196_c7_43ef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1196_c7_43ef_cond,
t8_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue,
t8_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse,
t8_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef
result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef
result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef
result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef
result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef
result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_cond,
result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c
BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_left,
BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_right,
BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_return_output);

-- n8_MUX_uxn_opcodes_h_l1199_c7_28f4
n8_MUX_uxn_opcodes_h_l1199_c7_28f4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1199_c7_28f4_cond,
n8_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue,
n8_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse,
n8_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4
result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4
result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4
result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_cond,
result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe
sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_ins,
sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_x,
sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_y,
sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1205_c21_4630
BIN_OP_EQ_uxn_opcodes_h_l1205_c21_4630 : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1205_c21_4630_left,
BIN_OP_EQ_uxn_opcodes_h_l1205_c21_4630_right,
BIN_OP_EQ_uxn_opcodes_h_l1205_c21_4630_return_output);

-- MUX_uxn_opcodes_h_l1205_c21_c121
MUX_uxn_opcodes_h_l1205_c21_c121 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1205_c21_c121_cond,
MUX_uxn_opcodes_h_l1205_c21_c121_iftrue,
MUX_uxn_opcodes_h_l1205_c21_c121_iffalse,
MUX_uxn_opcodes_h_l1205_c21_c121_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1207_c11_acd0
BIN_OP_EQ_uxn_opcodes_h_l1207_c11_acd0 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1207_c11_acd0_left,
BIN_OP_EQ_uxn_opcodes_h_l1207_c11_acd0_right,
BIN_OP_EQ_uxn_opcodes_h_l1207_c11_acd0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff
result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff
result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff
result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_return_output,
 n8_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output,
 t8_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_return_output,
 n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output,
 t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_return_output,
 n8_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output,
 t8_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_return_output,
 n8_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output,
 sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1205_c21_4630_return_output,
 MUX_uxn_opcodes_h_l1205_c21_c121_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1207_c11_acd0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1188_c2_a4da_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1188_c2_a4da_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1190_c3_a05a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1189_c3_7acb_uxn_opcodes_h_l1189_c3_7acb_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1194_c3_e431 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1196_c7_43ef_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1196_c7_43ef_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1199_c7_28f4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1204_c3_fe73 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1205_c21_c121_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1205_c21_c121_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1205_c21_c121_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_4630_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_4630_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_4630_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1205_c21_c121_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_acd0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_acd0_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_acd0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_3492_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_1014_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_40a3_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_2274_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1199_l1193_l1207_l1196_DUPLICATE_7bf1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1199_l1196_DUPLICATE_82c6_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1213_l1184_DUPLICATE_3f28_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_right := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_iffalse := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1205_c21_c121_iffalse := resize(to_unsigned(1, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1190_c3_a05a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1190_c3_a05a;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_acd0_right := to_unsigned(4, 3);
     VAR_MUX_uxn_opcodes_h_l1205_c21_c121_iftrue := resize(to_unsigned(0, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1194_c3_e431 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1194_c3_e431;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1204_c3_fe73 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1204_c3_fe73;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_acd0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_4630_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_4630_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_3492 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_3492_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1207_c11_acd0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1207_c11_acd0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_acd0_left;
     BIN_OP_EQ_uxn_opcodes_h_l1207_c11_acd0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_acd0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_acd0_return_output := BIN_OP_EQ_uxn_opcodes_h_l1207_c11_acd0_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1199_l1193_l1207_l1196_DUPLICATE_7bf1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1199_l1193_l1207_l1196_DUPLICATE_7bf1_return_output := result.is_opc_done;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_40a3 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_40a3_return_output := result.sp_relative_shift;

     -- sp_relative_shift[uxn_opcodes_h_l1202_c30_11fe] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_ins;
     sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_x;
     sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_return_output := sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1199_c11_f09c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_2274 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_2274_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1188_c6_a30b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1193_c11_c6fc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_left;
     BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_return_output := BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1196_c11_4891] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_left;
     BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_return_output := BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1205_c21_4630] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1205_c21_4630_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_4630_left;
     BIN_OP_EQ_uxn_opcodes_h_l1205_c21_4630_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_4630_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_4630_return_output := BIN_OP_EQ_uxn_opcodes_h_l1205_c21_4630_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_1014 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_1014_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1199_l1196_DUPLICATE_82c6 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1199_l1196_DUPLICATE_82c6_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1188_c2_a4da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1188_c2_a4da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_a30b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_c6fc_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1196_c7_43ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1196_c7_43ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_4891_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1199_c7_28f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_f09c_return_output;
     VAR_MUX_uxn_opcodes_h_l1205_c21_c121_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_4630_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_acd0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_acd0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_acd0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_40a3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_40a3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_40a3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_40a3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1199_l1193_l1207_l1196_DUPLICATE_7bf1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1199_l1193_l1207_l1196_DUPLICATE_7bf1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1199_l1193_l1207_l1196_DUPLICATE_7bf1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1199_l1193_l1207_l1196_DUPLICATE_7bf1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_1014_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_1014_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_1014_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_1014_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_3492_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_3492_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_3492_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1188_l1193_l1207_l1196_DUPLICATE_3492_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1199_l1196_DUPLICATE_82c6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1199_l1196_DUPLICATE_82c6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_2274_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_2274_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_2274_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1188_l1199_l1193_l1196_DUPLICATE_2274_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_11fe_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1199_c7_28f4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output;

     -- t8_MUX[uxn_opcodes_h_l1196_c7_43ef] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1196_c7_43ef_cond <= VAR_t8_MUX_uxn_opcodes_h_l1196_c7_43ef_cond;
     t8_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue;
     t8_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output := t8_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1207_c7_46ff] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1188_c1_1dc7] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1207_c7_46ff] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1207_c7_46ff] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_return_output;

     -- n8_MUX[uxn_opcodes_h_l1199_c7_28f4] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1199_c7_28f4_cond <= VAR_n8_MUX_uxn_opcodes_h_l1199_c7_28f4_cond;
     n8_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue;
     n8_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output := n8_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1199_c7_28f4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output;

     -- MUX[uxn_opcodes_h_l1205_c21_c121] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1205_c21_c121_cond <= VAR_MUX_uxn_opcodes_h_l1205_c21_c121_cond;
     MUX_uxn_opcodes_h_l1205_c21_c121_iftrue <= VAR_MUX_uxn_opcodes_h_l1205_c21_c121_iftrue;
     MUX_uxn_opcodes_h_l1205_c21_c121_iffalse <= VAR_MUX_uxn_opcodes_h_l1205_c21_c121_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1205_c21_c121_return_output := MUX_uxn_opcodes_h_l1205_c21_c121_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue := VAR_MUX_uxn_opcodes_h_l1205_c21_c121_return_output;
     VAR_printf_uxn_opcodes_h_l1189_c3_7acb_uxn_opcodes_h_l1189_c3_7acb_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_1dc7_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_46ff_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_46ff_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_46ff_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1199_c7_28f4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output;

     -- t8_MUX[uxn_opcodes_h_l1193_c7_cbcd] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond <= VAR_t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond;
     t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue;
     t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output := t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output;

     -- n8_MUX[uxn_opcodes_h_l1196_c7_43ef] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1196_c7_43ef_cond <= VAR_n8_MUX_uxn_opcodes_h_l1196_c7_43ef_cond;
     n8_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue;
     n8_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output := n8_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1199_c7_28f4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output := result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1196_c7_43ef] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1199_c7_28f4] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1196_c7_43ef] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output;

     -- printf_uxn_opcodes_h_l1189_c3_7acb[uxn_opcodes_h_l1189_c3_7acb] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1189_c3_7acb_uxn_opcodes_h_l1189_c3_7acb_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1189_c3_7acb_uxn_opcodes_h_l1189_c3_7acb_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1199_c7_28f4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_28f4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1196_c7_43ef] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1196_c7_43ef] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1193_c7_cbcd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output;

     -- t8_MUX[uxn_opcodes_h_l1188_c2_a4da] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1188_c2_a4da_cond <= VAR_t8_MUX_uxn_opcodes_h_l1188_c2_a4da_cond;
     t8_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue;
     t8_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output := t8_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1193_c7_cbcd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1196_c7_43ef] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output;

     -- n8_MUX[uxn_opcodes_h_l1193_c7_cbcd] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond <= VAR_n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond;
     n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue;
     n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output := n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1196_c7_43ef] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output := result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_43ef_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1188_c2_a4da] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1193_c7_cbcd] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output;

     -- n8_MUX[uxn_opcodes_h_l1188_c2_a4da] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1188_c2_a4da_cond <= VAR_n8_MUX_uxn_opcodes_h_l1188_c2_a4da_cond;
     n8_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue;
     n8_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output := n8_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1193_c7_cbcd] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1193_c7_cbcd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1193_c7_cbcd] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output := result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1188_c2_a4da] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_cbcd_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1188_c2_a4da] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1188_c2_a4da] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output := result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1188_c2_a4da] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1188_c2_a4da] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1213_l1184_DUPLICATE_3f28 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1213_l1184_DUPLICATE_3f28_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5b93(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_a4da_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1213_l1184_DUPLICATE_3f28_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1213_l1184_DUPLICATE_3f28_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
