-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 55
entity ldr_0CLK_a6885b22 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldr_0CLK_a6885b22;
architecture arch of ldr_0CLK_a6885b22 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1689_c6_bfde]
signal BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1689_c1_5951]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1689_c2_813f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_return_output : signed(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1689_c2_813f]
signal result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1689_c2_813f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1689_c2_813f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1689_c2_813f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1689_c2_813f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1689_c2_813f]
signal result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1689_c2_813f]
signal tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1689_c2_813f]
signal t8_MUX_uxn_opcodes_h_l1689_c2_813f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1689_c2_813f_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1690_c3_c5e5[uxn_opcodes_h_l1690_c3_c5e5]
signal printf_uxn_opcodes_h_l1690_c3_c5e5_uxn_opcodes_h_l1690_c3_c5e5_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1694_c11_52c8]
signal BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1694_c7_18db]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_return_output : signed(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1694_c7_18db]
signal result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1694_c7_18db]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1694_c7_18db]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1694_c7_18db]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1694_c7_18db]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1694_c7_18db]
signal result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1694_c7_18db]
signal tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1694_c7_18db]
signal t8_MUX_uxn_opcodes_h_l1694_c7_18db_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1694_c7_18db_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1697_c11_5d28]
signal BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1697_c7_37e7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output : signed(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1697_c7_37e7]
signal result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1697_c7_37e7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1697_c7_37e7]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1697_c7_37e7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1697_c7_37e7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1697_c7_37e7]
signal result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1697_c7_37e7]
signal tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1697_c7_37e7]
signal t8_MUX_uxn_opcodes_h_l1697_c7_37e7_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1700_c30_72d4]
signal sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_return_output : signed(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1701_c22_98d1]
signal BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_98d1_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_98d1_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_98d1_return_output : signed(17 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1703_c11_6442]
signal BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1703_c7_d096]
signal result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1703_c7_d096]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1703_c7_d096]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1703_c7_d096]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1703_c7_d096]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1703_c7_d096]
signal result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1703_c7_d096]
signal tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_return_output : unsigned(7 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1705_c22_2f53]
signal BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_2f53_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_2f53_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_2f53_return_output : signed(17 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1707_c11_fd4e]
signal BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1707_c7_885e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1707_c7_885e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1707_c7_885e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1707_c7_885e]
signal result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1707_c7_885e]
signal tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1713_c11_91e0]
signal BIN_OP_EQ_uxn_opcodes_h_l1713_c11_91e0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1713_c11_91e0_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1713_c11_91e0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1713_c7_6536]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1713_c7_6536]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_return_output : unsigned(0 downto 0);

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_1a88( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.u16_value := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_sp_shift := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.u8_value := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde
BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_left,
BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_right,
BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f
result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_cond,
result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f
result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f
result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f
result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f
result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1689_c2_813f
tmp8_MUX_uxn_opcodes_h_l1689_c2_813f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_cond,
tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue,
tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse,
tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_return_output);

-- t8_MUX_uxn_opcodes_h_l1689_c2_813f
t8_MUX_uxn_opcodes_h_l1689_c2_813f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1689_c2_813f_cond,
t8_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue,
t8_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse,
t8_MUX_uxn_opcodes_h_l1689_c2_813f_return_output);

-- printf_uxn_opcodes_h_l1690_c3_c5e5_uxn_opcodes_h_l1690_c3_c5e5
printf_uxn_opcodes_h_l1690_c3_c5e5_uxn_opcodes_h_l1690_c3_c5e5 : entity work.printf_uxn_opcodes_h_l1690_c3_c5e5_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1690_c3_c5e5_uxn_opcodes_h_l1690_c3_c5e5_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8
BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_left,
BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_right,
BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db
result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db
result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_cond,
result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db
result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db
result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db
result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db
result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_cond,
result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1694_c7_18db
tmp8_MUX_uxn_opcodes_h_l1694_c7_18db : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_cond,
tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue,
tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse,
tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_return_output);

-- t8_MUX_uxn_opcodes_h_l1694_c7_18db
t8_MUX_uxn_opcodes_h_l1694_c7_18db : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1694_c7_18db_cond,
t8_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue,
t8_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse,
t8_MUX_uxn_opcodes_h_l1694_c7_18db_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28
BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_left,
BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_right,
BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7
result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7
result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_cond,
result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7
result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7
result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7
result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7
result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_cond,
result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7
tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_cond,
tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue,
tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse,
tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output);

-- t8_MUX_uxn_opcodes_h_l1697_c7_37e7
t8_MUX_uxn_opcodes_h_l1697_c7_37e7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1697_c7_37e7_cond,
t8_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue,
t8_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse,
t8_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4
sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_ins,
sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_x,
sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_y,
sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_98d1
BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_98d1 : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_98d1_left,
BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_98d1_right,
BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_98d1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442
BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_left,
BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_right,
BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096
result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_cond,
result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096
result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096
result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096
result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096
result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_cond,
result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1703_c7_d096
tmp8_MUX_uxn_opcodes_h_l1703_c7_d096 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_cond,
tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue,
tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse,
tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_2f53
BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_2f53 : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_2f53_left,
BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_2f53_right,
BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_2f53_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e
BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e_left,
BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e_right,
BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e
result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e
result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e
result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_cond,
result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1707_c7_885e
tmp8_MUX_uxn_opcodes_h_l1707_c7_885e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_cond,
tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue,
tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse,
tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1713_c11_91e0
BIN_OP_EQ_uxn_opcodes_h_l1713_c11_91e0 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1713_c11_91e0_left,
BIN_OP_EQ_uxn_opcodes_h_l1713_c11_91e0_right,
BIN_OP_EQ_uxn_opcodes_h_l1713_c11_91e0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536
result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536
result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_return_output,
 tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_return_output,
 t8_MUX_uxn_opcodes_h_l1689_c2_813f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_return_output,
 tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_return_output,
 t8_MUX_uxn_opcodes_h_l1694_c7_18db_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output,
 tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output,
 t8_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output,
 sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_98d1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_return_output,
 tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_2f53_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_return_output,
 tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1713_c11_91e0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_iffalse : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1691_c3_9032 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1694_c7_18db_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1689_c2_813f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1689_c2_813f_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1690_c3_c5e5_uxn_opcodes_h_l1690_c3_c5e5_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1695_c3_2834 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1694_c7_18db_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l1701_c3_7e14 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1697_c7_37e7_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_98d1_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l1701_c27_4a7a_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_98d1_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_98d1_return_output : signed(17 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l1705_c3_cf61 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_2f53_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l1705_c27_bee6_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_2f53_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_2f53_return_output : signed(17 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1710_c3_fc3f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1713_c11_91e0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1713_c11_91e0_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1713_c11_91e0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1694_l1697_l1689_DUPLICATE_d2ec_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1694_l1689_l1703_DUPLICATE_02c4_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1694_l1689_l1703_DUPLICATE_141d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1703_l1697_l1694_l1689_l1713_DUPLICATE_fb64_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1707_l1703_l1697_l1694_l1689_DUPLICATE_e28d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1707_l1703_l1697_l1694_l1713_DUPLICATE_466f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1707_l1697_l1703_DUPLICATE_a797_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1a88_uxn_opcodes_h_l1685_l1718_DUPLICATE_7554_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1710_c3_fc3f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1710_c3_fc3f;
     VAR_sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1691_c3_9032 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1691_c3_9032;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1713_c11_91e0_right := to_unsigned(4, 3);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1695_c3_2834 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1695_c3_2834;
     VAR_sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_ins := VAR_ins;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_98d1_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_2f53_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1713_c11_91e0_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse := tmp8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1694_c11_52c8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_left;
     BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_return_output := BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1707_l1703_l1697_l1694_l1689_DUPLICATE_e28d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1707_l1703_l1697_l1694_l1689_DUPLICATE_e28d_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1703_c11_6442] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_left;
     BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_return_output := BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1700_c30_72d4] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_ins;
     sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_x;
     sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_return_output := sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1713_c11_91e0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1713_c11_91e0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1713_c11_91e0_left;
     BIN_OP_EQ_uxn_opcodes_h_l1713_c11_91e0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1713_c11_91e0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1713_c11_91e0_return_output := BIN_OP_EQ_uxn_opcodes_h_l1713_c11_91e0_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1694_l1689_l1703_DUPLICATE_02c4 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1694_l1689_l1703_DUPLICATE_02c4_return_output := result.u16_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1707_c11_fd4e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1707_l1703_l1697_l1694_l1713_DUPLICATE_466f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1707_l1703_l1697_l1694_l1713_DUPLICATE_466f_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1697_c11_5d28] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_left;
     BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_return_output := BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1689_c6_bfde] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_left;
     BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_return_output := BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1707_l1697_l1703_DUPLICATE_a797 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1707_l1697_l1703_DUPLICATE_a797_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1703_l1697_l1694_l1689_l1713_DUPLICATE_fb64 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1703_l1697_l1694_l1689_l1713_DUPLICATE_fb64_return_output := result.is_stack_write;

     -- CAST_TO_int8_t[uxn_opcodes_h_l1705_c27_bee6] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l1705_c27_bee6_return_output := CAST_TO_int8_t_uint8_t(
     t8);

     -- CAST_TO_int8_t[uxn_opcodes_h_l1701_c27_4a7a] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l1701_c27_4a7a_return_output := CAST_TO_int8_t_uint8_t(
     VAR_previous_stack_read);

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1694_l1697_l1689_DUPLICATE_d2ec LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1694_l1697_l1689_DUPLICATE_d2ec_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1694_l1689_l1703_DUPLICATE_141d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1694_l1689_l1703_DUPLICATE_141d_return_output := result.is_sp_shift;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1689_c2_813f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_bfde_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1694_c7_18db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_52c8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1697_c7_37e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_5d28_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_6442_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_fd4e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1713_c11_91e0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1713_c11_91e0_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_98d1_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l1701_c27_4a7a_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_2f53_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l1705_c27_bee6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1694_l1697_l1689_DUPLICATE_d2ec_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1694_l1697_l1689_DUPLICATE_d2ec_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1694_l1697_l1689_DUPLICATE_d2ec_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1694_l1689_l1703_DUPLICATE_02c4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1694_l1689_l1703_DUPLICATE_02c4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1694_l1689_l1703_DUPLICATE_02c4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1707_l1703_l1697_l1694_l1713_DUPLICATE_466f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1707_l1703_l1697_l1694_l1713_DUPLICATE_466f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1707_l1703_l1697_l1694_l1713_DUPLICATE_466f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1707_l1703_l1697_l1694_l1713_DUPLICATE_466f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1707_l1703_l1697_l1694_l1713_DUPLICATE_466f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1694_l1689_l1703_DUPLICATE_141d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1694_l1689_l1703_DUPLICATE_141d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1694_l1689_l1703_DUPLICATE_141d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1703_l1697_l1694_l1689_l1713_DUPLICATE_fb64_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1703_l1697_l1694_l1689_l1713_DUPLICATE_fb64_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1703_l1697_l1694_l1689_l1713_DUPLICATE_fb64_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1703_l1697_l1694_l1689_l1713_DUPLICATE_fb64_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1703_l1697_l1694_l1689_l1713_DUPLICATE_fb64_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1707_l1697_l1703_DUPLICATE_a797_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1707_l1697_l1703_DUPLICATE_a797_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1707_l1697_l1703_DUPLICATE_a797_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1707_l1703_l1697_l1694_l1689_DUPLICATE_e28d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1707_l1703_l1697_l1694_l1689_DUPLICATE_e28d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1707_l1703_l1697_l1694_l1689_DUPLICATE_e28d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1707_l1703_l1697_l1694_l1689_DUPLICATE_e28d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1707_l1703_l1697_l1694_l1689_DUPLICATE_e28d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1700_c30_72d4_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1713_c7_6536] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1707_c7_885e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1697_c7_37e7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1713_c7_6536] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1705_c22_2f53] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_2f53_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_2f53_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_2f53_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_2f53_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_2f53_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_2f53_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1703_c7_d096] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_return_output;

     -- t8_MUX[uxn_opcodes_h_l1697_c7_37e7] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1697_c7_37e7_cond <= VAR_t8_MUX_uxn_opcodes_h_l1697_c7_37e7_cond;
     t8_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue;
     t8_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output := t8_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1707_c7_885e] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_cond;
     tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_return_output := tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1707_c7_885e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_return_output := result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1701_c22_98d1] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_98d1_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_98d1_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_98d1_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_98d1_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_98d1_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_98d1_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1689_c1_5951] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_return_output;

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l1701_c3_7e14 := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_98d1_return_output)),16);
     VAR_result_u16_value_uxn_opcodes_h_l1705_c3_cf61 := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_2f53_return_output)),16);
     VAR_printf_uxn_opcodes_h_l1690_c3_c5e5_uxn_opcodes_h_l1690_c3_c5e5_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_5951_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_6536_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_d096_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_6536_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_885e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1707_c7_885e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1707_c7_885e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue := VAR_result_u16_value_uxn_opcodes_h_l1701_c3_7e14;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue := VAR_result_u16_value_uxn_opcodes_h_l1705_c3_cf61;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1697_c7_37e7] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output;

     -- printf_uxn_opcodes_h_l1690_c3_c5e5[uxn_opcodes_h_l1690_c3_c5e5] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1690_c3_c5e5_uxn_opcodes_h_l1690_c3_c5e5_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1690_c3_c5e5_uxn_opcodes_h_l1690_c3_c5e5_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- tmp8_MUX[uxn_opcodes_h_l1703_c7_d096] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_cond;
     tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_return_output := tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1707_c7_885e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1694_c7_18db] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1703_c7_d096] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_return_output := result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_return_output;

     -- t8_MUX[uxn_opcodes_h_l1694_c7_18db] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1694_c7_18db_cond <= VAR_t8_MUX_uxn_opcodes_h_l1694_c7_18db_cond;
     t8_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue;
     t8_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1694_c7_18db_return_output := t8_MUX_uxn_opcodes_h_l1694_c7_18db_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1703_c7_d096] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_return_output := result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1703_c7_d096] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1707_c7_885e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_885e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_885e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_18db_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_d096_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_d096_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_d096_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1694_c7_18db_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1703_c7_d096_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1703_c7_d096] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1697_c7_37e7] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_cond;
     tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output := tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1694_c7_18db] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1703_c7_d096] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1689_c2_813f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1697_c7_37e7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output := result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output;

     -- t8_MUX[uxn_opcodes_h_l1689_c2_813f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1689_c2_813f_cond <= VAR_t8_MUX_uxn_opcodes_h_l1689_c2_813f_cond;
     t8_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue;
     t8_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1689_c2_813f_return_output := t8_MUX_uxn_opcodes_h_l1689_c2_813f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1697_c7_37e7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1697_c7_37e7] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output := result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_d096_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_18db_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_d096_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1689_c2_813f_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1694_c7_18db] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_return_output := result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1694_c7_18db] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1697_c7_37e7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1689_c2_813f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1694_c7_18db] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_return_output := result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1694_c7_18db] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_cond;
     tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_return_output := tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1697_c7_37e7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_37e7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_18db_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c7_18db_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c7_18db_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1694_c7_18db_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1694_c7_18db] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1694_c7_18db] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1689_c2_813f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1689_c2_813f] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_cond;
     tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_return_output := tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1689_c2_813f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1689_c2_813f] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_return_output := result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_18db_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_18db_return_output;
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1689_c2_813f_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1689_c2_813f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1689_c2_813f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_1a88_uxn_opcodes_h_l1685_l1718_DUPLICATE_7554 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1a88_uxn_opcodes_h_l1685_l1718_DUPLICATE_7554_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_1a88(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_813f_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1689_c2_813f_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_813f_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_813f_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_813f_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_813f_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1689_c2_813f_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1a88_uxn_opcodes_h_l1685_l1718_DUPLICATE_7554_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1a88_uxn_opcodes_h_l1685_l1718_DUPLICATE_7554_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
