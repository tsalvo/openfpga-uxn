-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity stz_0CLK_bacf6a1d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end stz_0CLK_bacf6a1d;
architecture arch of stz_0CLK_bacf6a1d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1522_c6_e493]
signal BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1522_c2_6696]
signal n8_MUX_uxn_opcodes_h_l1522_c2_6696_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1522_c2_6696]
signal result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1522_c2_6696]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1522_c2_6696]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1522_c2_6696]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1522_c2_6696]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1522_c2_6696]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1522_c2_6696]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1522_c2_6696]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1522_c2_6696]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1522_c2_6696]
signal result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1522_c2_6696]
signal t8_MUX_uxn_opcodes_h_l1522_c2_6696_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1535_c11_9a31]
signal BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1535_c7_5ad2]
signal n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1535_c7_5ad2]
signal result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1535_c7_5ad2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1535_c7_5ad2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1535_c7_5ad2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1535_c7_5ad2]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1535_c7_5ad2]
signal result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1535_c7_5ad2]
signal t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1538_c11_109b]
signal BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1538_c7_dad7]
signal n8_MUX_uxn_opcodes_h_l1538_c7_dad7_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1538_c7_dad7]
signal result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1538_c7_dad7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1538_c7_dad7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1538_c7_dad7]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1538_c7_dad7]
signal result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1538_c7_dad7]
signal t8_MUX_uxn_opcodes_h_l1538_c7_dad7_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1541_c11_99db]
signal BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1541_c7_9a3d]
signal n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1541_c7_9a3d]
signal result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1541_c7_9a3d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1541_c7_9a3d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1541_c7_9a3d]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1541_c7_9a3d]
signal result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1543_c30_662f]
signal sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_return_output : signed(3 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_a906( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u16_value := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.stack_address_sp_offset := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_vram_write := ref_toks_8;
      base.is_pc_updated := ref_toks_9;
      base.u8_value := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493
BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_left,
BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_right,
BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_return_output);

-- n8_MUX_uxn_opcodes_h_l1522_c2_6696
n8_MUX_uxn_opcodes_h_l1522_c2_6696 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1522_c2_6696_cond,
n8_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue,
n8_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse,
n8_MUX_uxn_opcodes_h_l1522_c2_6696_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696
result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_cond,
result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696
result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696
result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696
result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696
result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696
result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696
result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696
result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_cond,
result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_return_output);

-- t8_MUX_uxn_opcodes_h_l1522_c2_6696
t8_MUX_uxn_opcodes_h_l1522_c2_6696 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1522_c2_6696_cond,
t8_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue,
t8_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse,
t8_MUX_uxn_opcodes_h_l1522_c2_6696_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31
BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_left,
BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_right,
BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_return_output);

-- n8_MUX_uxn_opcodes_h_l1535_c7_5ad2
n8_MUX_uxn_opcodes_h_l1535_c7_5ad2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond,
n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue,
n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse,
n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2
result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond,
result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2
result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2
result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2
result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2
result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond,
result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output);

-- t8_MUX_uxn_opcodes_h_l1535_c7_5ad2
t8_MUX_uxn_opcodes_h_l1535_c7_5ad2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond,
t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue,
t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse,
t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b
BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_left,
BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_right,
BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_return_output);

-- n8_MUX_uxn_opcodes_h_l1538_c7_dad7
n8_MUX_uxn_opcodes_h_l1538_c7_dad7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1538_c7_dad7_cond,
n8_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue,
n8_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse,
n8_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7
result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_cond,
result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7
result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7
result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7
result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7
result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_cond,
result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output);

-- t8_MUX_uxn_opcodes_h_l1538_c7_dad7
t8_MUX_uxn_opcodes_h_l1538_c7_dad7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1538_c7_dad7_cond,
t8_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue,
t8_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse,
t8_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db
BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db_left,
BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db_right,
BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db_return_output);

-- n8_MUX_uxn_opcodes_h_l1541_c7_9a3d
n8_MUX_uxn_opcodes_h_l1541_c7_9a3d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond,
n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue,
n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse,
n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d
result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond,
result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d
result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d
result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d
result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d
result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond,
result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1543_c30_662f
sp_relative_shift_uxn_opcodes_h_l1543_c30_662f : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_ins,
sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_x,
sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_y,
sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_return_output,
 n8_MUX_uxn_opcodes_h_l1522_c2_6696_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_return_output,
 t8_MUX_uxn_opcodes_h_l1522_c2_6696_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_return_output,
 n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output,
 t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_return_output,
 n8_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output,
 t8_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db_return_output,
 n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output,
 sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1522_c2_6696_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1532_c3_d4f5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1527_c3_a329 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1522_c2_6696_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1522_c2_6696_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1536_c3_8540 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1535_c7_5ad2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1538_c7_dad7_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1538_c7_dad7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1545_c22_f6b9_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1522_l1541_l1535_l1538_DUPLICATE_dadc_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1522_l1541_l1535_l1538_DUPLICATE_e9b5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1541_l1535_l1538_DUPLICATE_3fca_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1541_l1535_l1538_DUPLICATE_16b8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1541_l1535_l1538_DUPLICATE_e5e7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a906_uxn_opcodes_h_l1550_l1518_DUPLICATE_7803_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1527_c3_a329 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1527_c3_a329;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_y := resize(to_signed(-2, 3), 4);
     VAR_sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1532_c3_d4f5 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1532_c3_d4f5;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1536_c3_8540 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1536_c3_8540;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_right := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse := t8;
     -- CAST_TO_uint16_t[uxn_opcodes_h_l1545_c22_f6b9] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1545_c22_f6b9_return_output := CAST_TO_uint16_t_uint8_t(
     t8);

     -- BIN_OP_EQ[uxn_opcodes_h_l1538_c11_109b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1543_c30_662f] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_ins;
     sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_x;
     sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_return_output := sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1522_c2_6696] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1522_c2_6696_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1522_l1541_l1535_l1538_DUPLICATE_e9b5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1522_l1541_l1535_l1538_DUPLICATE_e9b5_return_output := result.u8_value;

     -- result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d[uxn_opcodes_h_l1522_c2_6696] LATENCY=0
     VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1522_c2_6696_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1541_l1535_l1538_DUPLICATE_e5e7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1541_l1535_l1538_DUPLICATE_e5e7_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1541_l1535_l1538_DUPLICATE_16b8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1541_l1535_l1538_DUPLICATE_16b8_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1522_l1541_l1535_l1538_DUPLICATE_dadc LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1522_l1541_l1535_l1538_DUPLICATE_dadc_return_output := result.u16_value;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1522_c2_6696] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1522_c2_6696_return_output := result.is_pc_updated;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1535_c7_5ad2] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1535_c7_5ad2_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1535_c11_9a31] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_left;
     BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_return_output := BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1541_c11_99db] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db_left;
     BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db_return_output := BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1541_l1535_l1538_DUPLICATE_3fca LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1541_l1535_l1538_DUPLICATE_3fca_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1522_c6_e493] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_left;
     BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_return_output := BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1522_c2_6696] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1522_c2_6696_return_output := result.is_stack_index_flipped;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1522_c2_6696_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1522_c2_6696_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1522_c6_e493_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1535_c11_9a31_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1538_c7_dad7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1538_c7_dad7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_109b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_99db_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1545_c22_f6b9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1541_l1535_l1538_DUPLICATE_3fca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1541_l1535_l1538_DUPLICATE_3fca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1541_l1535_l1538_DUPLICATE_3fca_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1522_l1541_l1535_l1538_DUPLICATE_dadc_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1522_l1541_l1535_l1538_DUPLICATE_dadc_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1522_l1541_l1535_l1538_DUPLICATE_dadc_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1522_l1541_l1535_l1538_DUPLICATE_dadc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1541_l1535_l1538_DUPLICATE_16b8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1541_l1535_l1538_DUPLICATE_16b8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1541_l1535_l1538_DUPLICATE_16b8_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1541_l1535_l1538_DUPLICATE_e5e7_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1541_l1535_l1538_DUPLICATE_e5e7_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1541_l1535_l1538_DUPLICATE_e5e7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1522_l1541_l1535_l1538_DUPLICATE_e9b5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1522_l1541_l1535_l1538_DUPLICATE_e9b5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1522_l1541_l1535_l1538_DUPLICATE_e9b5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1522_l1541_l1535_l1538_DUPLICATE_e9b5_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1522_c2_6696_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1522_c2_6696_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse := VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1522_c2_6696_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1522_c2_6696_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1535_c7_5ad2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1543_c30_662f_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1522_c2_6696] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_return_output;

     -- t8_MUX[uxn_opcodes_h_l1538_c7_dad7] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1538_c7_dad7_cond <= VAR_t8_MUX_uxn_opcodes_h_l1538_c7_dad7_cond;
     t8_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue;
     t8_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output := t8_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1541_c7_9a3d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1541_c7_9a3d] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output := result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1522_c2_6696] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1541_c7_9a3d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1541_c7_9a3d] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1522_c2_6696] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_return_output;

     -- n8_MUX[uxn_opcodes_h_l1541_c7_9a3d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond <= VAR_n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond;
     n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue;
     n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output := n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1522_c2_6696] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1541_c7_9a3d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output := result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1535_c7_5ad2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_9a3d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1538_c7_dad7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1538_c7_dad7] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1522_c2_6696] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1538_c7_dad7] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output := result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1538_c7_dad7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output := result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output;

     -- n8_MUX[uxn_opcodes_h_l1538_c7_dad7] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1538_c7_dad7_cond <= VAR_n8_MUX_uxn_opcodes_h_l1538_c7_dad7_cond;
     n8_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue;
     n8_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output := n8_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1538_c7_dad7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output;

     -- t8_MUX[uxn_opcodes_h_l1535_c7_5ad2] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond <= VAR_t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond;
     t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue;
     t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output := t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1538_c7_dad7_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1535_c7_5ad2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output;

     -- n8_MUX[uxn_opcodes_h_l1535_c7_5ad2] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond <= VAR_n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond;
     n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue;
     n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output := n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1535_c7_5ad2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output := result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output;

     -- t8_MUX[uxn_opcodes_h_l1522_c2_6696] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1522_c2_6696_cond <= VAR_t8_MUX_uxn_opcodes_h_l1522_c2_6696_cond;
     t8_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue;
     t8_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1522_c2_6696_return_output := t8_MUX_uxn_opcodes_h_l1522_c2_6696_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1535_c7_5ad2] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1535_c7_5ad2] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output := result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1535_c7_5ad2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1535_c7_5ad2_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1522_c2_6696_return_output;
     -- result_is_ram_write_MUX[uxn_opcodes_h_l1522_c2_6696] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_return_output;

     -- n8_MUX[uxn_opcodes_h_l1522_c2_6696] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1522_c2_6696_cond <= VAR_n8_MUX_uxn_opcodes_h_l1522_c2_6696_cond;
     n8_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue;
     n8_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1522_c2_6696_return_output := n8_MUX_uxn_opcodes_h_l1522_c2_6696_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1522_c2_6696] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_return_output := result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1522_c2_6696] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1522_c2_6696] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1522_c2_6696] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_return_output := result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1522_c2_6696_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a906_uxn_opcodes_h_l1550_l1518_DUPLICATE_7803 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a906_uxn_opcodes_h_l1550_l1518_DUPLICATE_7803_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a906(
     result,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1522_c2_6696_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1522_c2_6696_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1522_c2_6696_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1522_c2_6696_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1522_c2_6696_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1522_c2_6696_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1522_c2_6696_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1522_c2_6696_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1522_c2_6696_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1522_c2_6696_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a906_uxn_opcodes_h_l1550_l1518_DUPLICATE_7803_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a906_uxn_opcodes_h_l1550_l1518_DUPLICATE_7803_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
