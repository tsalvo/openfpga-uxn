-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity jsr_0CLK_6d7675a8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jsr_0CLK_6d7675a8;
architecture arch of jsr_0CLK_6d7675a8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l722_c6_ab48]
signal BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l722_c2_2ec1]
signal result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l722_c2_2ec1]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l722_c2_2ec1]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l722_c2_2ec1]
signal result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l722_c2_2ec1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l722_c2_2ec1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l722_c2_2ec1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l722_c2_2ec1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l722_c2_2ec1]
signal t8_MUX_uxn_opcodes_h_l722_c2_2ec1_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l729_c11_7d90]
signal BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l729_c7_75c6]
signal result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l729_c7_75c6]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l729_c7_75c6]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l729_c7_75c6]
signal result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l729_c7_75c6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l729_c7_75c6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l729_c7_75c6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l729_c7_75c6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l729_c7_75c6]
signal t8_MUX_uxn_opcodes_h_l729_c7_75c6_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l729_c7_75c6_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l732_c30_7c2d]
signal sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l734_c11_dc21]
signal BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l734_c7_8f3e]
signal result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l734_c7_8f3e]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l734_c7_8f3e]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l734_c7_8f3e]
signal result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l734_c7_8f3e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l734_c7_8f3e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l734_c7_8f3e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l734_c7_8f3e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l734_c7_8f3e]
signal t8_MUX_uxn_opcodes_h_l734_c7_8f3e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l742_c11_f22f]
signal BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l742_c7_1c13]
signal result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l742_c7_1c13]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l742_c7_1c13]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l742_c7_1c13]
signal result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l742_c7_1c13]
signal result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l742_c7_1c13]
signal result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l742_c7_1c13]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l742_c7_1c13]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_return_output : unsigned(3 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l745_c31_a7d1]
signal CONST_SR_8_uxn_opcodes_h_l745_c31_a7d1_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l745_c31_a7d1_return_output : unsigned(15 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l747_c22_7c57]
signal BIN_OP_PLUS_uxn_opcodes_h_l747_c22_7c57_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l747_c22_7c57_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l747_c22_7c57_return_output : signed(17 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l749_c11_eddd]
signal BIN_OP_EQ_uxn_opcodes_h_l749_c11_eddd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l749_c11_eddd_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l749_c11_eddd_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l749_c7_9a35]
signal result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l749_c7_9a35]
signal result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l749_c7_9a35]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l749_c7_9a35]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_return_output : unsigned(0 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_a30a( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.is_pc_updated := ref_toks_3;
      base.u16_value := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.is_opc_done := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48
BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_left,
BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_right,
BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1
result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_cond,
result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1
result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1
result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_cond,
result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1
result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1
result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1
result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output);

-- t8_MUX_uxn_opcodes_h_l722_c2_2ec1
t8_MUX_uxn_opcodes_h_l722_c2_2ec1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l722_c2_2ec1_cond,
t8_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue,
t8_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse,
t8_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90
BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_left,
BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_right,
BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6
result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_cond,
result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6
result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6
result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_cond,
result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6
result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6
result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6
result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_return_output);

-- t8_MUX_uxn_opcodes_h_l729_c7_75c6
t8_MUX_uxn_opcodes_h_l729_c7_75c6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l729_c7_75c6_cond,
t8_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue,
t8_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse,
t8_MUX_uxn_opcodes_h_l729_c7_75c6_return_output);

-- sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d
sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_ins,
sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_x,
sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_y,
sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21
BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_left,
BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_right,
BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e
result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_cond,
result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e
result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e
result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_cond,
result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e
result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e
result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e
result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output);

-- t8_MUX_uxn_opcodes_h_l734_c7_8f3e
t8_MUX_uxn_opcodes_h_l734_c7_8f3e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l734_c7_8f3e_cond,
t8_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue,
t8_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse,
t8_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f
BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_left,
BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_right,
BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13
result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_cond,
result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13
result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13
result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_cond,
result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13
result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13
result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13
result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_return_output);

-- CONST_SR_8_uxn_opcodes_h_l745_c31_a7d1
CONST_SR_8_uxn_opcodes_h_l745_c31_a7d1 : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l745_c31_a7d1_x,
CONST_SR_8_uxn_opcodes_h_l745_c31_a7d1_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l747_c22_7c57
BIN_OP_PLUS_uxn_opcodes_h_l747_c22_7c57 : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l747_c22_7c57_left,
BIN_OP_PLUS_uxn_opcodes_h_l747_c22_7c57_right,
BIN_OP_PLUS_uxn_opcodes_h_l747_c22_7c57_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l749_c11_eddd
BIN_OP_EQ_uxn_opcodes_h_l749_c11_eddd : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l749_c11_eddd_left,
BIN_OP_EQ_uxn_opcodes_h_l749_c11_eddd_right,
BIN_OP_EQ_uxn_opcodes_h_l749_c11_eddd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35
result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35
result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35
result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output,
 t8_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_return_output,
 t8_MUX_uxn_opcodes_h_l729_c7_75c6_return_output,
 sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output,
 t8_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_return_output,
 CONST_SR_8_uxn_opcodes_h_l745_c31_a7d1_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l747_c22_7c57_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l749_c11_eddd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l726_c3_7158 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l729_c7_75c6_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l722_c2_2ec1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l730_c3_6d26 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l729_c7_75c6_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l737_c3_94e0 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l739_c3_9a0c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l734_c7_8f3e_cond : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l740_c21_8960_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l747_c3_acf5 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l743_c3_fd78 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l744_c3_14ea : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l742_c7_1c13_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l745_c31_a7d1_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l745_c31_a7d1_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l745_c21_ac4c_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l747_c22_7c57_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l747_c27_c9c8_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l747_c22_7c57_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l747_c22_7c57_return_output : signed(17 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_eddd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_eddd_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_eddd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l729_l722_l742_DUPLICATE_3ba4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l729_l749_l722_l742_DUPLICATE_c245_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l729_l749_l734_l722_DUPLICATE_057d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l729_l734_l722_l742_DUPLICATE_999f_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l729_l749_l722_l742_DUPLICATE_5a95_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l722_l742_DUPLICATE_f5a3_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l729_l749_l734_l742_DUPLICATE_8ccd_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a30a_uxn_opcodes_h_l756_l718_DUPLICATE_42bf_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l730_c3_6d26 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l730_c3_6d26;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_eddd_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l744_c3_14ea := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l744_c3_14ea;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l726_c3_7158 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l726_c3_7158;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l739_c3_9a0c := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l739_c3_9a0c;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_y := resize(to_signed(-1, 2), 4);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l737_c3_94e0 := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l737_c3_94e0;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_right := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l743_c3_fd78 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l743_c3_fd78;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_ins := VAR_ins;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l747_c22_7c57_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_CONST_SR_8_uxn_opcodes_h_l745_c31_a7d1_x := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_eddd_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse := t8;
     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l729_l722_l742_DUPLICATE_3ba4 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l729_l722_l742_DUPLICATE_3ba4_return_output := result.u8_value;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l729_l734_l722_l742_DUPLICATE_999f LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l729_l734_l722_l742_DUPLICATE_999f_return_output := result.u16_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l729_l749_l734_l722_DUPLICATE_057d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l729_l749_l734_l722_DUPLICATE_057d_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l722_c6_ab48] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_left;
     BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_return_output := BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l734_c11_dc21] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_left;
     BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_return_output := BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l729_l749_l722_l742_DUPLICATE_c245 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l729_l749_l722_l742_DUPLICATE_c245_return_output := result.is_stack_index_flipped;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l742_c7_1c13] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l742_c7_1c13_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l729_c11_7d90] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_left;
     BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_return_output := BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_return_output;

     -- CAST_TO_int8_t[uxn_opcodes_h_l747_c27_c9c8] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l747_c27_c9c8_return_output := CAST_TO_int8_t_uint8_t(
     t8);

     -- CONST_SR_8[uxn_opcodes_h_l745_c31_a7d1] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l745_c31_a7d1_x <= VAR_CONST_SR_8_uxn_opcodes_h_l745_c31_a7d1_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l745_c31_a7d1_return_output := CONST_SR_8_uxn_opcodes_h_l745_c31_a7d1_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l732_c30_7c2d] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_ins;
     sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_x <= VAR_sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_x;
     sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_y <= VAR_sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_return_output := sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l729_l749_l722_l742_DUPLICATE_5a95 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l729_l749_l722_l742_DUPLICATE_5a95_return_output := result.is_stack_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l722_l742_DUPLICATE_f5a3 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l722_l742_DUPLICATE_f5a3_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l749_c11_eddd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l749_c11_eddd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_eddd_left;
     BIN_OP_EQ_uxn_opcodes_h_l749_c11_eddd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_eddd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_eddd_return_output := BIN_OP_EQ_uxn_opcodes_h_l749_c11_eddd_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l742_c11_f22f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_left;
     BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_return_output := BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l740_c21_8960] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l740_c21_8960_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_pc);

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l729_l749_l734_l742_DUPLICATE_8ccd LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l729_l749_l734_l742_DUPLICATE_8ccd_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l722_c2_2ec1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l722_c6_ab48_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l729_c7_75c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l729_c11_7d90_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l734_c7_8f3e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l734_c11_dc21_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l742_c11_f22f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_eddd_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_eddd_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_eddd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_eddd_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l747_c22_7c57_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l747_c27_c9c8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l740_c21_8960_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l722_l742_DUPLICATE_f5a3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l722_l742_DUPLICATE_f5a3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l729_l734_l722_l742_DUPLICATE_999f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l729_l734_l722_l742_DUPLICATE_999f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l729_l734_l722_l742_DUPLICATE_999f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l729_l734_l722_l742_DUPLICATE_999f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l729_l749_l734_l742_DUPLICATE_8ccd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l729_l749_l734_l742_DUPLICATE_8ccd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l729_l749_l734_l742_DUPLICATE_8ccd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l729_l749_l734_l742_DUPLICATE_8ccd_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l729_l749_l734_l722_DUPLICATE_057d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l729_l749_l734_l722_DUPLICATE_057d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l729_l749_l734_l722_DUPLICATE_057d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l729_l749_l734_l722_DUPLICATE_057d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l729_l749_l722_l742_DUPLICATE_c245_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l729_l749_l722_l742_DUPLICATE_c245_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l729_l749_l722_l742_DUPLICATE_c245_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l729_l749_l722_l742_DUPLICATE_c245_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l729_l749_l722_l742_DUPLICATE_5a95_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l729_l749_l722_l742_DUPLICATE_5a95_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l729_l749_l722_l742_DUPLICATE_5a95_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l729_l749_l722_l742_DUPLICATE_5a95_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l729_l722_l742_DUPLICATE_3ba4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l729_l722_l742_DUPLICATE_3ba4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l729_l722_l742_DUPLICATE_3ba4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l742_c7_1c13_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l732_c30_7c2d_return_output;
     -- t8_MUX[uxn_opcodes_h_l734_c7_8f3e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l734_c7_8f3e_cond <= VAR_t8_MUX_uxn_opcodes_h_l734_c7_8f3e_cond;
     t8_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue;
     t8_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output := t8_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l747_c22_7c57] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l747_c22_7c57_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l747_c22_7c57_left;
     BIN_OP_PLUS_uxn_opcodes_h_l747_c22_7c57_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l747_c22_7c57_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l747_c22_7c57_return_output := BIN_OP_PLUS_uxn_opcodes_h_l747_c22_7c57_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l749_c7_9a35] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l749_c7_9a35] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l749_c7_9a35] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l742_c7_1c13] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l742_c7_1c13] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l749_c7_9a35] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l745_c21_ac4c] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l745_c21_ac4c_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l745_c31_a7d1_return_output);

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l747_c3_acf5 := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l747_c22_7c57_return_output)),16);
     VAR_result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l745_c21_ac4c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_9a35_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_9a35_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_9a35_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_9a35_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l742_c7_1c13_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l742_c7_1c13_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse := VAR_t8_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue := VAR_result_u16_value_uxn_opcodes_h_l747_c3_acf5;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l742_c7_1c13] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l742_c7_1c13] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_cond;
     result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_return_output := result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l742_c7_1c13] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l742_c7_1c13] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l734_c7_8f3e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l734_c7_8f3e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l742_c7_1c13] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_cond;
     result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_return_output := result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_return_output;

     -- t8_MUX[uxn_opcodes_h_l729_c7_75c6] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l729_c7_75c6_cond <= VAR_t8_MUX_uxn_opcodes_h_l729_c7_75c6_cond;
     t8_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue;
     t8_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l729_c7_75c6_return_output := t8_MUX_uxn_opcodes_h_l729_c7_75c6_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l742_c7_1c13] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l742_c7_1c13_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l742_c7_1c13_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l742_c7_1c13_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l742_c7_1c13_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l742_c7_1c13_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l742_c7_1c13_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse := VAR_t8_MUX_uxn_opcodes_h_l729_c7_75c6_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l734_c7_8f3e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output := result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l734_c7_8f3e] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l734_c7_8f3e] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_cond;
     result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output := result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l729_c7_75c6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l729_c7_75c6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_return_output;

     -- t8_MUX[uxn_opcodes_h_l722_c2_2ec1] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l722_c2_2ec1_cond <= VAR_t8_MUX_uxn_opcodes_h_l722_c2_2ec1_cond;
     t8_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue;
     t8_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output := t8_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l734_c7_8f3e] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l734_c7_8f3e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l734_c7_8f3e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l729_c7_75c6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l729_c7_75c6_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l734_c7_8f3e_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l729_c7_75c6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l729_c7_75c6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_return_output := result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l729_c7_75c6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l722_c2_2ec1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l729_c7_75c6] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_cond;
     result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_return_output := result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l729_c7_75c6] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l729_c7_75c6] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l722_c2_2ec1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l729_c7_75c6_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l729_c7_75c6_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l729_c7_75c6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l729_c7_75c6_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l729_c7_75c6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l729_c7_75c6_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l722_c2_2ec1] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_cond;
     result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output := result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l722_c2_2ec1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l722_c2_2ec1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l722_c2_2ec1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output := result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l722_c2_2ec1] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l722_c2_2ec1] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a30a_uxn_opcodes_h_l756_l718_DUPLICATE_42bf LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a30a_uxn_opcodes_h_l756_l718_DUPLICATE_42bf_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a30a(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l722_c2_2ec1_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a30a_uxn_opcodes_h_l756_l718_DUPLICATE_42bf_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a30a_uxn_opcodes_h_l756_l718_DUPLICATE_42bf_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
