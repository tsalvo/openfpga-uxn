-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity ovr_0CLK_61914e8d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ovr_0CLK_61914e8d;
architecture arch of ovr_0CLK_61914e8d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l297_c6_3b4b]
signal BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l297_c2_e657]
signal n8_MUX_uxn_opcodes_h_l297_c2_e657_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l297_c2_e657_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l297_c2_e657_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l297_c2_e657_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l297_c2_e657]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l297_c2_e657]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l297_c2_e657]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l297_c2_e657]
signal result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l297_c2_e657]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l297_c2_e657]
signal result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l297_c2_e657]
signal result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l297_c2_e657]
signal result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l297_c2_e657]
signal result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l297_c2_e657]
signal t8_MUX_uxn_opcodes_h_l297_c2_e657_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l297_c2_e657_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l297_c2_e657_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l297_c2_e657_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l310_c11_77c6]
signal BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l310_c7_248d]
signal n8_MUX_uxn_opcodes_h_l310_c7_248d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l310_c7_248d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l310_c7_248d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l310_c7_248d_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l310_c7_248d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l310_c7_248d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l310_c7_248d]
signal result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l310_c7_248d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l310_c7_248d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l310_c7_248d]
signal t8_MUX_uxn_opcodes_h_l310_c7_248d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l310_c7_248d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l310_c7_248d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l310_c7_248d_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l313_c11_7295]
signal BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l313_c7_affd]
signal n8_MUX_uxn_opcodes_h_l313_c7_affd_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l313_c7_affd_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l313_c7_affd_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l313_c7_affd_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l313_c7_affd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l313_c7_affd]
signal result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l313_c7_affd]
signal result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l313_c7_affd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l313_c7_affd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l313_c7_affd]
signal t8_MUX_uxn_opcodes_h_l313_c7_affd_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l313_c7_affd_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l313_c7_affd_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l313_c7_affd_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l315_c30_cca4]
signal sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l320_c11_259f]
signal BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l320_c7_be36]
signal n8_MUX_uxn_opcodes_h_l320_c7_be36_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l320_c7_be36_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l320_c7_be36_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l320_c7_be36_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l320_c7_be36]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l320_c7_be36]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l320_c7_be36]
signal result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l320_c7_be36]
signal result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l326_c11_a6ad]
signal BIN_OP_EQ_uxn_opcodes_h_l326_c11_a6ad_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l326_c11_a6ad_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l326_c11_a6ad_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l326_c7_5cdb]
signal result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l326_c7_5cdb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l326_c7_5cdb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8b52( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_opc_done := ref_toks_6;
      base.is_ram_write := ref_toks_7;
      base.is_vram_write := ref_toks_8;
      base.u8_value := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b
BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_left,
BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_right,
BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_return_output);

-- n8_MUX_uxn_opcodes_h_l297_c2_e657
n8_MUX_uxn_opcodes_h_l297_c2_e657 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l297_c2_e657_cond,
n8_MUX_uxn_opcodes_h_l297_c2_e657_iftrue,
n8_MUX_uxn_opcodes_h_l297_c2_e657_iffalse,
n8_MUX_uxn_opcodes_h_l297_c2_e657_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657
result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_cond,
result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_return_output);

-- t8_MUX_uxn_opcodes_h_l297_c2_e657
t8_MUX_uxn_opcodes_h_l297_c2_e657 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l297_c2_e657_cond,
t8_MUX_uxn_opcodes_h_l297_c2_e657_iftrue,
t8_MUX_uxn_opcodes_h_l297_c2_e657_iffalse,
t8_MUX_uxn_opcodes_h_l297_c2_e657_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6
BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_left,
BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_right,
BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_return_output);

-- n8_MUX_uxn_opcodes_h_l310_c7_248d
n8_MUX_uxn_opcodes_h_l310_c7_248d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l310_c7_248d_cond,
n8_MUX_uxn_opcodes_h_l310_c7_248d_iftrue,
n8_MUX_uxn_opcodes_h_l310_c7_248d_iffalse,
n8_MUX_uxn_opcodes_h_l310_c7_248d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d
result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_cond,
result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_return_output);

-- t8_MUX_uxn_opcodes_h_l310_c7_248d
t8_MUX_uxn_opcodes_h_l310_c7_248d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l310_c7_248d_cond,
t8_MUX_uxn_opcodes_h_l310_c7_248d_iftrue,
t8_MUX_uxn_opcodes_h_l310_c7_248d_iffalse,
t8_MUX_uxn_opcodes_h_l310_c7_248d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295
BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_left,
BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_right,
BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_return_output);

-- n8_MUX_uxn_opcodes_h_l313_c7_affd
n8_MUX_uxn_opcodes_h_l313_c7_affd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l313_c7_affd_cond,
n8_MUX_uxn_opcodes_h_l313_c7_affd_iftrue,
n8_MUX_uxn_opcodes_h_l313_c7_affd_iffalse,
n8_MUX_uxn_opcodes_h_l313_c7_affd_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd
result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_cond,
result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_return_output);

-- t8_MUX_uxn_opcodes_h_l313_c7_affd
t8_MUX_uxn_opcodes_h_l313_c7_affd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l313_c7_affd_cond,
t8_MUX_uxn_opcodes_h_l313_c7_affd_iftrue,
t8_MUX_uxn_opcodes_h_l313_c7_affd_iffalse,
t8_MUX_uxn_opcodes_h_l313_c7_affd_return_output);

-- sp_relative_shift_uxn_opcodes_h_l315_c30_cca4
sp_relative_shift_uxn_opcodes_h_l315_c30_cca4 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_ins,
sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_x,
sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_y,
sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f
BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f_left,
BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f_right,
BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f_return_output);

-- n8_MUX_uxn_opcodes_h_l320_c7_be36
n8_MUX_uxn_opcodes_h_l320_c7_be36 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l320_c7_be36_cond,
n8_MUX_uxn_opcodes_h_l320_c7_be36_iftrue,
n8_MUX_uxn_opcodes_h_l320_c7_be36_iffalse,
n8_MUX_uxn_opcodes_h_l320_c7_be36_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36
result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_cond,
result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l326_c11_a6ad
BIN_OP_EQ_uxn_opcodes_h_l326_c11_a6ad : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l326_c11_a6ad_left,
BIN_OP_EQ_uxn_opcodes_h_l326_c11_a6ad_right,
BIN_OP_EQ_uxn_opcodes_h_l326_c11_a6ad_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb
result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_cond,
result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_return_output,
 n8_MUX_uxn_opcodes_h_l297_c2_e657_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_return_output,
 t8_MUX_uxn_opcodes_h_l297_c2_e657_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_return_output,
 n8_MUX_uxn_opcodes_h_l310_c7_248d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_return_output,
 t8_MUX_uxn_opcodes_h_l310_c7_248d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_return_output,
 n8_MUX_uxn_opcodes_h_l313_c7_affd_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_return_output,
 t8_MUX_uxn_opcodes_h_l313_c7_affd_return_output,
 sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f_return_output,
 n8_MUX_uxn_opcodes_h_l320_c7_be36_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l326_c11_a6ad_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l297_c2_e657_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l297_c2_e657_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l310_c7_248d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l297_c2_e657_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l297_c2_e657_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l302_c3_0510 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l297_c2_e657_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l297_c2_e657_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l307_c3_8fdc : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l297_c2_e657_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l297_c2_e657_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l297_c2_e657_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l297_c2_e657_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l310_c7_248d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l297_c2_e657_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l297_c2_e657_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l310_c7_248d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l310_c7_248d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l313_c7_affd_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l310_c7_248d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l311_c3_2878 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l310_c7_248d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l310_c7_248d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l313_c7_affd_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l310_c7_248d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l313_c7_affd_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l313_c7_affd_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l320_c7_be36_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l313_c7_affd_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l317_c3_87da : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l313_c7_affd_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l313_c7_affd_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l313_c7_affd_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l320_c7_be36_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l320_c7_be36_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l320_c7_be36_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l323_c3_e6ec : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l322_c3_5162 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_a6ad_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_a6ad_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_a6ad_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l327_c3_75c4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l326_c7_5cdb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l326_l297_l310_DUPLICATE_389d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l320_l310_DUPLICATE_2197_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l313_l310_DUPLICATE_5fdf_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l313_l326_l320_l310_DUPLICATE_66aa_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l293_l332_DUPLICATE_000c_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_a6ad_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l302_c3_0510 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l302_c3_0510;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l327_c3_75c4 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l327_c3_75c4;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l322_c3_5162 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l322_c3_5162;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l317_c3_87da := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l317_c3_87da;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l323_c3_e6ec := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l323_c3_e6ec;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l307_c3_8fdc := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l307_c3_8fdc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l311_c3_2878 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l311_c3_2878;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l297_c2_e657_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l310_c7_248d_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l313_c7_affd_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l320_c7_be36_iffalse := n8;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_iftrue := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_a6ad_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l320_c7_be36_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l313_c7_affd_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l297_c2_e657_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l310_c7_248d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l313_c7_affd_iffalse := t8;
     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l326_l297_l310_DUPLICATE_389d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l326_l297_l310_DUPLICATE_389d_return_output := result.u8_value;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l297_c2_e657] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l297_c2_e657_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l313_c11_7295] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_left;
     BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_return_output := BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l326_c7_5cdb] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l326_c7_5cdb_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l326_c11_a6ad] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l326_c11_a6ad_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_a6ad_left;
     BIN_OP_EQ_uxn_opcodes_h_l326_c11_a6ad_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_a6ad_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_a6ad_return_output := BIN_OP_EQ_uxn_opcodes_h_l326_c11_a6ad_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l297_c6_3b4b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_left;
     BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_return_output := BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l315_c30_cca4] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_ins;
     sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_x <= VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_x;
     sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_y <= VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_return_output := sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l320_l310_DUPLICATE_2197 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l320_l310_DUPLICATE_2197_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l313_l310_DUPLICATE_5fdf LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l313_l310_DUPLICATE_5fdf_return_output := result.is_stack_write;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l297_c2_e657] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l297_c2_e657_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l310_c11_77c6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_left;
     BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_return_output := BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l313_l326_l320_l310_DUPLICATE_66aa LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l313_l326_l320_l310_DUPLICATE_66aa_return_output := result.is_opc_done;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l297_c2_e657] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l297_c2_e657_return_output := result.is_ram_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l297_c2_e657] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l297_c2_e657_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l320_c11_259f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f_left;
     BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f_return_output := BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l297_c2_e657_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l297_c2_e657_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_3b4b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l310_c7_248d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l310_c7_248d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_77c6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l313_c7_affd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l313_c7_affd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_7295_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l320_c7_be36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_259f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_a6ad_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_a6ad_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_a6ad_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l320_l310_DUPLICATE_2197_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l320_l310_DUPLICATE_2197_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l313_l326_l320_l310_DUPLICATE_66aa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l313_l326_l320_l310_DUPLICATE_66aa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l313_l326_l320_l310_DUPLICATE_66aa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l313_l326_l320_l310_DUPLICATE_66aa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l313_l310_DUPLICATE_5fdf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l313_l310_DUPLICATE_5fdf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l326_l297_l310_DUPLICATE_389d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l326_l297_l310_DUPLICATE_389d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l326_l297_l310_DUPLICATE_389d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l297_c2_e657_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l297_c2_e657_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l297_c2_e657_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l297_c2_e657_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l326_c7_5cdb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_cca4_return_output;
     -- t8_MUX[uxn_opcodes_h_l313_c7_affd] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l313_c7_affd_cond <= VAR_t8_MUX_uxn_opcodes_h_l313_c7_affd_cond;
     t8_MUX_uxn_opcodes_h_l313_c7_affd_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l313_c7_affd_iftrue;
     t8_MUX_uxn_opcodes_h_l313_c7_affd_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l313_c7_affd_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l313_c7_affd_return_output := t8_MUX_uxn_opcodes_h_l313_c7_affd_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l297_c2_e657] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l297_c2_e657] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l326_c7_5cdb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l297_c2_e657] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l326_c7_5cdb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l320_c7_be36] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l313_c7_affd] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l297_c2_e657] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l326_c7_5cdb] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_cond;
     result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_return_output := result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_return_output;

     -- n8_MUX[uxn_opcodes_h_l320_c7_be36] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l320_c7_be36_cond <= VAR_n8_MUX_uxn_opcodes_h_l320_c7_be36_cond;
     n8_MUX_uxn_opcodes_h_l320_c7_be36_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l320_c7_be36_iftrue;
     n8_MUX_uxn_opcodes_h_l320_c7_be36_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l320_c7_be36_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l320_c7_be36_return_output := n8_MUX_uxn_opcodes_h_l320_c7_be36_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l313_c7_affd_iffalse := VAR_n8_MUX_uxn_opcodes_h_l320_c7_be36_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_5cdb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_affd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_be36_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_5cdb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_5cdb_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l310_c7_248d_iffalse := VAR_t8_MUX_uxn_opcodes_h_l313_c7_affd_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l310_c7_248d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l320_c7_be36] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_return_output;

     -- t8_MUX[uxn_opcodes_h_l310_c7_248d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l310_c7_248d_cond <= VAR_t8_MUX_uxn_opcodes_h_l310_c7_248d_cond;
     t8_MUX_uxn_opcodes_h_l310_c7_248d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l310_c7_248d_iftrue;
     t8_MUX_uxn_opcodes_h_l310_c7_248d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l310_c7_248d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l310_c7_248d_return_output := t8_MUX_uxn_opcodes_h_l310_c7_248d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l313_c7_affd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l320_c7_be36] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_cond;
     result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_return_output := result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l320_c7_be36] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_return_output;

     -- n8_MUX[uxn_opcodes_h_l313_c7_affd] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l313_c7_affd_cond <= VAR_n8_MUX_uxn_opcodes_h_l313_c7_affd_cond;
     n8_MUX_uxn_opcodes_h_l313_c7_affd_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l313_c7_affd_iftrue;
     n8_MUX_uxn_opcodes_h_l313_c7_affd_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l313_c7_affd_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l313_c7_affd_return_output := n8_MUX_uxn_opcodes_h_l313_c7_affd_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l310_c7_248d_iffalse := VAR_n8_MUX_uxn_opcodes_h_l313_c7_affd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_be36_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_248d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_affd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_be36_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_be36_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l297_c2_e657_iffalse := VAR_t8_MUX_uxn_opcodes_h_l310_c7_248d_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l313_c7_affd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_return_output;

     -- t8_MUX[uxn_opcodes_h_l297_c2_e657] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l297_c2_e657_cond <= VAR_t8_MUX_uxn_opcodes_h_l297_c2_e657_cond;
     t8_MUX_uxn_opcodes_h_l297_c2_e657_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l297_c2_e657_iftrue;
     t8_MUX_uxn_opcodes_h_l297_c2_e657_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l297_c2_e657_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l297_c2_e657_return_output := t8_MUX_uxn_opcodes_h_l297_c2_e657_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l310_c7_248d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l313_c7_affd] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_cond;
     result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_return_output := result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_return_output;

     -- n8_MUX[uxn_opcodes_h_l310_c7_248d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l310_c7_248d_cond <= VAR_n8_MUX_uxn_opcodes_h_l310_c7_248d_cond;
     n8_MUX_uxn_opcodes_h_l310_c7_248d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l310_c7_248d_iftrue;
     n8_MUX_uxn_opcodes_h_l310_c7_248d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l310_c7_248d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l310_c7_248d_return_output := n8_MUX_uxn_opcodes_h_l310_c7_248d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l313_c7_affd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l297_c2_e657] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l297_c2_e657_iffalse := VAR_n8_MUX_uxn_opcodes_h_l310_c7_248d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_affd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_248d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_affd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_affd_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l297_c2_e657_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l297_c2_e657] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l310_c7_248d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_return_output;

     -- n8_MUX[uxn_opcodes_h_l297_c2_e657] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l297_c2_e657_cond <= VAR_n8_MUX_uxn_opcodes_h_l297_c2_e657_cond;
     n8_MUX_uxn_opcodes_h_l297_c2_e657_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l297_c2_e657_iftrue;
     n8_MUX_uxn_opcodes_h_l297_c2_e657_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l297_c2_e657_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l297_c2_e657_return_output := n8_MUX_uxn_opcodes_h_l297_c2_e657_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l310_c7_248d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_return_output := result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l310_c7_248d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l297_c2_e657_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_248d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_248d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_248d_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l297_c2_e657] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l297_c2_e657] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l297_c2_e657] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_cond;
     result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_return_output := result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l293_l332_DUPLICATE_000c LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l293_l332_DUPLICATE_000c_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8b52(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_e657_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_e657_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_e657_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_e657_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_e657_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_e657_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_e657_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_e657_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_e657_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l293_l332_DUPLICATE_000c_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l293_l332_DUPLICATE_000c_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
