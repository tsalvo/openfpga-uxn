-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 41
entity str1_0CLK_85d5529e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end str1_0CLK_85d5529e;
architecture arch of str1_0CLK_85d5529e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1705_c6_5480]
signal BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1705_c2_94ff]
signal n8_MUX_uxn_opcodes_h_l1705_c2_94ff_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1705_c2_94ff]
signal t8_MUX_uxn_opcodes_h_l1705_c2_94ff_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1705_c2_94ff]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1705_c2_94ff]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1705_c2_94ff]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1705_c2_94ff]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1705_c2_94ff]
signal result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1705_c2_94ff]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1705_c2_94ff]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1705_c2_94ff]
signal result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1705_c2_94ff]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1705_c2_94ff]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1718_c11_d06f]
signal BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1718_c7_6812]
signal n8_MUX_uxn_opcodes_h_l1718_c7_6812_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1718_c7_6812_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1718_c7_6812]
signal t8_MUX_uxn_opcodes_h_l1718_c7_6812_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1718_c7_6812_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1718_c7_6812]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_return_output : unsigned(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1718_c7_6812]
signal result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1718_c7_6812]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1718_c7_6812]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1718_c7_6812]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1718_c7_6812]
signal result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1721_c11_02a9]
signal BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1721_c7_4d3a]
signal n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1721_c7_4d3a]
signal t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1721_c7_4d3a]
signal result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1721_c7_4d3a]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1721_c7_4d3a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1721_c7_4d3a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1721_c7_4d3a]
signal result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1724_c11_62ad]
signal BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1724_c7_17dd]
signal n8_MUX_uxn_opcodes_h_l1724_c7_17dd_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1724_c7_17dd]
signal result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1724_c7_17dd]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1724_c7_17dd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1724_c7_17dd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1724_c7_17dd]
signal result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1726_c30_9499]
signal sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_return_output : signed(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1728_c22_95b2]
signal BIN_OP_PLUS_uxn_opcodes_h_l1728_c22_95b2_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1728_c22_95b2_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1728_c22_95b2_return_output : signed(17 downto 0);

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_vram_write := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;
      base.u16_value := ref_toks_8;
      base.is_pc_updated := ref_toks_9;
      base.is_opc_done := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480
BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_left,
BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_right,
BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_return_output);

-- n8_MUX_uxn_opcodes_h_l1705_c2_94ff
n8_MUX_uxn_opcodes_h_l1705_c2_94ff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1705_c2_94ff_cond,
n8_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue,
n8_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse,
n8_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output);

-- t8_MUX_uxn_opcodes_h_l1705_c2_94ff
t8_MUX_uxn_opcodes_h_l1705_c2_94ff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1705_c2_94ff_cond,
t8_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue,
t8_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse,
t8_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff
result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff
result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff
result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff
result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff
result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_cond,
result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff
result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_cond,
result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff
result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff
result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f
BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_left,
BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_right,
BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_return_output);

-- n8_MUX_uxn_opcodes_h_l1718_c7_6812
n8_MUX_uxn_opcodes_h_l1718_c7_6812 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1718_c7_6812_cond,
n8_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue,
n8_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse,
n8_MUX_uxn_opcodes_h_l1718_c7_6812_return_output);

-- t8_MUX_uxn_opcodes_h_l1718_c7_6812
t8_MUX_uxn_opcodes_h_l1718_c7_6812 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1718_c7_6812_cond,
t8_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue,
t8_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse,
t8_MUX_uxn_opcodes_h_l1718_c7_6812_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812
result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_cond,
result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812
result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812
result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812
result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812
result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_cond,
result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9
BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_left,
BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_right,
BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_return_output);

-- n8_MUX_uxn_opcodes_h_l1721_c7_4d3a
n8_MUX_uxn_opcodes_h_l1721_c7_4d3a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond,
n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue,
n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse,
n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output);

-- t8_MUX_uxn_opcodes_h_l1721_c7_4d3a
t8_MUX_uxn_opcodes_h_l1721_c7_4d3a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond,
t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue,
t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse,
t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a
result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond,
result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a
result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a
result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a
result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a
result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond,
result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad
BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad_left,
BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad_right,
BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad_return_output);

-- n8_MUX_uxn_opcodes_h_l1724_c7_17dd
n8_MUX_uxn_opcodes_h_l1724_c7_17dd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1724_c7_17dd_cond,
n8_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue,
n8_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse,
n8_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd
result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_cond,
result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd
result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd
result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd
result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd
result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_cond,
result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1726_c30_9499
sp_relative_shift_uxn_opcodes_h_l1726_c30_9499 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_ins,
sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_x,
sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_y,
sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1728_c22_95b2
BIN_OP_PLUS_uxn_opcodes_h_l1728_c22_95b2 : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1728_c22_95b2_left,
BIN_OP_PLUS_uxn_opcodes_h_l1728_c22_95b2_right,
BIN_OP_PLUS_uxn_opcodes_h_l1728_c22_95b2_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_return_output,
 n8_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output,
 t8_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_return_output,
 n8_MUX_uxn_opcodes_h_l1718_c7_6812_return_output,
 t8_MUX_uxn_opcodes_h_l1718_c7_6812_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_return_output,
 n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output,
 t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad_return_output,
 n8_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output,
 sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1728_c22_95b2_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1718_c7_6812_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1705_c2_94ff_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1718_c7_6812_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1705_c2_94ff_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1710_c3_a761 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1715_c3_d100 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1718_c7_6812_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1718_c7_6812_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1719_c3_7eb7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1718_c7_6812_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1724_c7_17dd_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l1728_c3_191f : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1728_c22_95b2_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l1728_c27_c6c2_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1728_c22_95b2_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1728_c22_95b2_return_output : signed(17 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1718_l1721_l1705_l1724_DUPLICATE_66cf_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1718_l1721_l1705_l1724_DUPLICATE_3c85_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1718_l1721_l1724_DUPLICATE_d1e5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1718_l1721_l1724_DUPLICATE_24a5_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1718_l1721_l1724_DUPLICATE_aa7e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4_uxn_opcodes_h_l1733_l1701_DUPLICATE_09a9_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_y := resize(to_signed(-2, 3), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1719_c3_7eb7 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1719_c3_7eb7;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1710_c3_a761 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1710_c3_a761;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_right := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1715_c3_d100 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1715_c3_d100;
     VAR_sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse := n8;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1728_c22_95b2_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse := t8;
     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1718_l1721_l1705_l1724_DUPLICATE_3c85 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1718_l1721_l1705_l1724_DUPLICATE_3c85_return_output := result.u16_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1718_c11_d06f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1705_c2_94ff] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1705_c2_94ff_return_output := result.is_vram_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1705_c2_94ff] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1705_c2_94ff_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l1705_c6_5480] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_left;
     BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_return_output := BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1718_l1721_l1724_DUPLICATE_d1e5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1718_l1721_l1724_DUPLICATE_d1e5_return_output := result.is_ram_write;

     -- sp_relative_shift[uxn_opcodes_h_l1726_c30_9499] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_ins;
     sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_x;
     sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_return_output := sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1718_l1721_l1724_DUPLICATE_aa7e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1718_l1721_l1724_DUPLICATE_aa7e_return_output := result.is_opc_done;

     -- CAST_TO_int8_t[uxn_opcodes_h_l1728_c27_c6c2] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l1728_c27_c6c2_return_output := CAST_TO_int8_t_uint8_t(
     t8);

     -- result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d[uxn_opcodes_h_l1705_c2_94ff] LATENCY=0
     VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1705_c2_94ff_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1724_c11_62ad] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad_left;
     BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad_return_output := BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1718_l1721_l1724_DUPLICATE_24a5 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1718_l1721_l1724_DUPLICATE_24a5_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1721_c11_02a9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_left;
     BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_return_output := BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1718_c7_6812] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1718_c7_6812_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1718_l1721_l1705_l1724_DUPLICATE_66cf LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1718_l1721_l1705_l1724_DUPLICATE_66cf_return_output := result.u8_value;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1705_c2_94ff] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1705_c2_94ff_return_output := result.is_stack_index_flipped;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1705_c2_94ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1705_c2_94ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1705_c6_5480_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1718_c7_6812_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1718_c7_6812_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1718_c11_d06f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1721_c11_02a9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1724_c7_17dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1724_c11_62ad_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1728_c22_95b2_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l1728_c27_c6c2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1718_l1721_l1724_DUPLICATE_24a5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1718_l1721_l1724_DUPLICATE_24a5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1718_l1721_l1724_DUPLICATE_24a5_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1718_l1721_l1705_l1724_DUPLICATE_3c85_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1718_l1721_l1705_l1724_DUPLICATE_3c85_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1718_l1721_l1705_l1724_DUPLICATE_3c85_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1718_l1721_l1705_l1724_DUPLICATE_3c85_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1718_l1721_l1724_DUPLICATE_aa7e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1718_l1721_l1724_DUPLICATE_aa7e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1718_l1721_l1724_DUPLICATE_aa7e_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1718_l1721_l1724_DUPLICATE_d1e5_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1718_l1721_l1724_DUPLICATE_d1e5_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1718_l1721_l1724_DUPLICATE_d1e5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1718_l1721_l1705_l1724_DUPLICATE_66cf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1718_l1721_l1705_l1724_DUPLICATE_66cf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1718_l1721_l1705_l1724_DUPLICATE_66cf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1718_l1721_l1705_l1724_DUPLICATE_66cf_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1705_c2_94ff_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1705_c2_94ff_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse := VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1705_c2_94ff_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1705_c2_94ff_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1718_c7_6812_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1726_c30_9499_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1724_c7_17dd] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output := result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1728_c22_95b2] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1728_c22_95b2_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1728_c22_95b2_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1728_c22_95b2_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1728_c22_95b2_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1728_c22_95b2_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1728_c22_95b2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1705_c2_94ff] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1724_c7_17dd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1724_c7_17dd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1705_c2_94ff] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1705_c2_94ff] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1724_c7_17dd] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1718_c7_6812] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_return_output;

     -- n8_MUX[uxn_opcodes_h_l1724_c7_17dd] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1724_c7_17dd_cond <= VAR_n8_MUX_uxn_opcodes_h_l1724_c7_17dd_cond;
     n8_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue;
     n8_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output := n8_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1705_c2_94ff] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output;

     -- t8_MUX[uxn_opcodes_h_l1721_c7_4d3a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond <= VAR_t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond;
     t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue;
     t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output := t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output;

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l1728_c3_191f := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1728_c22_95b2_return_output)),16);
     VAR_n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1718_c7_6812_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue := VAR_result_u16_value_uxn_opcodes_h_l1728_c3_191f;
     -- n8_MUX[uxn_opcodes_h_l1721_c7_4d3a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond <= VAR_n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond;
     n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue;
     n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output := n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1721_c7_4d3a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output := result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1721_c7_4d3a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1721_c7_4d3a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1705_c2_94ff] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output;

     -- t8_MUX[uxn_opcodes_h_l1718_c7_6812] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1718_c7_6812_cond <= VAR_t8_MUX_uxn_opcodes_h_l1718_c7_6812_cond;
     t8_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue;
     t8_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1718_c7_6812_return_output := t8_MUX_uxn_opcodes_h_l1718_c7_6812_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1721_c7_4d3a] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1724_c7_17dd] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output := result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1724_c7_17dd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1718_c7_6812_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1718_c7_6812] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1718_c7_6812] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_return_output := result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_return_output;

     -- t8_MUX[uxn_opcodes_h_l1705_c2_94ff] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1705_c2_94ff_cond <= VAR_t8_MUX_uxn_opcodes_h_l1705_c2_94ff_cond;
     t8_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue;
     t8_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output := t8_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1721_c7_4d3a] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output := result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1718_c7_6812] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1718_c7_6812] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_return_output;

     -- n8_MUX[uxn_opcodes_h_l1718_c7_6812] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1718_c7_6812_cond <= VAR_n8_MUX_uxn_opcodes_h_l1718_c7_6812_cond;
     n8_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue;
     n8_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1718_c7_6812_return_output := n8_MUX_uxn_opcodes_h_l1718_c7_6812_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1718_c7_6812_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1718_c7_6812_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1718_c7_6812_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1718_c7_6812_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1721_c7_4d3a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1718_c7_6812_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l1718_c7_6812] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_return_output := result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1705_c2_94ff] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1705_c2_94ff] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output;

     -- n8_MUX[uxn_opcodes_h_l1705_c2_94ff] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1705_c2_94ff_cond <= VAR_n8_MUX_uxn_opcodes_h_l1705_c2_94ff_cond;
     n8_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue;
     n8_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output := n8_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1705_c2_94ff] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output := result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1705_c2_94ff] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1718_c7_6812_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l1705_c2_94ff] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output := result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4_uxn_opcodes_h_l1733_l1701_DUPLICATE_09a9 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4_uxn_opcodes_h_l1733_l1701_DUPLICATE_09a9_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1705_c2_94ff_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4_uxn_opcodes_h_l1733_l1701_DUPLICATE_09a9_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_dfe4_uxn_opcodes_h_l1733_l1701_DUPLICATE_09a9_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
