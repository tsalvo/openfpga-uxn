-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 46
entity div_0CLK_a35230ee is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end div_0CLK_a35230ee;
architecture arch of div_0CLK_a35230ee is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1953_c6_f299]
signal BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1953_c1_fcb0]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1953_c2_8dca]
signal t8_MUX_uxn_opcodes_h_l1953_c2_8dca_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1953_c2_8dca]
signal n8_MUX_uxn_opcodes_h_l1953_c2_8dca_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1953_c2_8dca]
signal result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1953_c2_8dca]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1953_c2_8dca]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1953_c2_8dca]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1953_c2_8dca]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1953_c2_8dca]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output : signed(3 downto 0);

-- printf_uxn_opcodes_h_l1954_c3_53b9[uxn_opcodes_h_l1954_c3_53b9]
signal printf_uxn_opcodes_h_l1954_c3_53b9_uxn_opcodes_h_l1954_c3_53b9_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1958_c11_6068]
signal BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1958_c7_c9d8]
signal t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1958_c7_c9d8]
signal n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1958_c7_c9d8]
signal result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1958_c7_c9d8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1958_c7_c9d8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1958_c7_c9d8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1958_c7_c9d8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1958_c7_c9d8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1961_c11_a553]
signal BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1961_c7_1b7a]
signal t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1961_c7_1b7a]
signal n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1961_c7_1b7a]
signal result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1961_c7_1b7a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1961_c7_1b7a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1961_c7_1b7a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1961_c7_1b7a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1961_c7_1b7a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1964_c11_3e14]
signal BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1964_c7_96da]
signal n8_MUX_uxn_opcodes_h_l1964_c7_96da_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1964_c7_96da_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1964_c7_96da]
signal result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1964_c7_96da]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1964_c7_96da]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1964_c7_96da]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1964_c7_96da]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1964_c7_96da]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_return_output : signed(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1967_c30_4d76]
signal sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1970_c21_a00d]
signal BIN_OP_EQ_uxn_opcodes_h_l1970_c21_a00d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1970_c21_a00d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1970_c21_a00d_return_output : unsigned(0 downto 0);

-- BIN_OP_DIV[uxn_opcodes_h_l1970_c35_bf62]
signal BIN_OP_DIV_uxn_opcodes_h_l1970_c35_bf62_left : unsigned(7 downto 0);
signal BIN_OP_DIV_uxn_opcodes_h_l1970_c35_bf62_right : unsigned(7 downto 0);
signal BIN_OP_DIV_uxn_opcodes_h_l1970_c35_bf62_return_output : unsigned(7 downto 0);

-- MUX[uxn_opcodes_h_l1970_c21_1af7]
signal MUX_uxn_opcodes_h_l1970_c21_1af7_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1970_c21_1af7_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1970_c21_1af7_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1970_c21_1af7_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1972_c11_374c]
signal BIN_OP_EQ_uxn_opcodes_h_l1972_c11_374c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1972_c11_374c_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1972_c11_374c_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1972_c7_9e83]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1972_c7_9e83]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1972_c7_9e83]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299
BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_left,
BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_right,
BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_return_output);

-- t8_MUX_uxn_opcodes_h_l1953_c2_8dca
t8_MUX_uxn_opcodes_h_l1953_c2_8dca : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1953_c2_8dca_cond,
t8_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue,
t8_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse,
t8_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output);

-- n8_MUX_uxn_opcodes_h_l1953_c2_8dca
n8_MUX_uxn_opcodes_h_l1953_c2_8dca : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1953_c2_8dca_cond,
n8_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue,
n8_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse,
n8_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca
result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_cond,
result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca
result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca
result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca
result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca
result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output);

-- printf_uxn_opcodes_h_l1954_c3_53b9_uxn_opcodes_h_l1954_c3_53b9
printf_uxn_opcodes_h_l1954_c3_53b9_uxn_opcodes_h_l1954_c3_53b9 : entity work.printf_uxn_opcodes_h_l1954_c3_53b9_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1954_c3_53b9_uxn_opcodes_h_l1954_c3_53b9_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068
BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_left,
BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_right,
BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_return_output);

-- t8_MUX_uxn_opcodes_h_l1958_c7_c9d8
t8_MUX_uxn_opcodes_h_l1958_c7_c9d8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond,
t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue,
t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse,
t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output);

-- n8_MUX_uxn_opcodes_h_l1958_c7_c9d8
n8_MUX_uxn_opcodes_h_l1958_c7_c9d8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond,
n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue,
n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse,
n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8
result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond,
result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8
result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8
result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8
result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8
result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553
BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_left,
BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_right,
BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_return_output);

-- t8_MUX_uxn_opcodes_h_l1961_c7_1b7a
t8_MUX_uxn_opcodes_h_l1961_c7_1b7a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond,
t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue,
t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse,
t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output);

-- n8_MUX_uxn_opcodes_h_l1961_c7_1b7a
n8_MUX_uxn_opcodes_h_l1961_c7_1b7a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond,
n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue,
n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse,
n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a
result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond,
result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a
result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a
result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a
result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a
result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14
BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_left,
BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_right,
BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_return_output);

-- n8_MUX_uxn_opcodes_h_l1964_c7_96da
n8_MUX_uxn_opcodes_h_l1964_c7_96da : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1964_c7_96da_cond,
n8_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue,
n8_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse,
n8_MUX_uxn_opcodes_h_l1964_c7_96da_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da
result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_cond,
result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da
result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da
result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da
result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da
result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76
sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_ins,
sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_x,
sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_y,
sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1970_c21_a00d
BIN_OP_EQ_uxn_opcodes_h_l1970_c21_a00d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1970_c21_a00d_left,
BIN_OP_EQ_uxn_opcodes_h_l1970_c21_a00d_right,
BIN_OP_EQ_uxn_opcodes_h_l1970_c21_a00d_return_output);

-- BIN_OP_DIV_uxn_opcodes_h_l1970_c35_bf62
BIN_OP_DIV_uxn_opcodes_h_l1970_c35_bf62 : entity work.BIN_OP_DIV_uint8_t_uint8_t_0CLK_a148083c port map (
BIN_OP_DIV_uxn_opcodes_h_l1970_c35_bf62_left,
BIN_OP_DIV_uxn_opcodes_h_l1970_c35_bf62_right,
BIN_OP_DIV_uxn_opcodes_h_l1970_c35_bf62_return_output);

-- MUX_uxn_opcodes_h_l1970_c21_1af7
MUX_uxn_opcodes_h_l1970_c21_1af7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1970_c21_1af7_cond,
MUX_uxn_opcodes_h_l1970_c21_1af7_iftrue,
MUX_uxn_opcodes_h_l1970_c21_1af7_iffalse,
MUX_uxn_opcodes_h_l1970_c21_1af7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1972_c11_374c
BIN_OP_EQ_uxn_opcodes_h_l1972_c11_374c : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1972_c11_374c_left,
BIN_OP_EQ_uxn_opcodes_h_l1972_c11_374c_right,
BIN_OP_EQ_uxn_opcodes_h_l1972_c11_374c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83
result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83
result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83
result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_return_output,
 t8_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output,
 n8_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_return_output,
 t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output,
 n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_return_output,
 t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output,
 n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_return_output,
 n8_MUX_uxn_opcodes_h_l1964_c7_96da_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_return_output,
 sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1970_c21_a00d_return_output,
 BIN_OP_DIV_uxn_opcodes_h_l1970_c35_bf62_return_output,
 MUX_uxn_opcodes_h_l1970_c21_1af7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1972_c11_374c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1953_c2_8dca_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1953_c2_8dca_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1955_c3_9fc5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1954_c3_53b9_uxn_opcodes_h_l1954_c3_53b9_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1959_c3_f12d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1964_c7_96da_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1964_c7_96da_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1969_c3_2858 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1970_c21_1af7_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1970_c21_1af7_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1970_c21_1af7_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c21_a00d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c21_a00d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c21_a00d_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l1970_c35_bf62_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l1970_c35_bf62_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l1970_c35_bf62_return_output : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1970_c21_1af7_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_374c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_374c_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_374c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1961_l1953_l1964_l1958_DUPLICATE_22d5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1961_l1953_l1958_l1972_DUPLICATE_21a0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1961_l1953_l1958_l1972_DUPLICATE_3e93_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1961_l1953_l1964_l1958_DUPLICATE_62fe_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1961_l1964_l1958_l1972_DUPLICATE_3cd0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1961_l1964_DUPLICATE_2fdb_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1978_l1949_DUPLICATE_1c81_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1969_c3_2858 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1969_c3_2858;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1959_c3_f12d := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1959_c3_f12d;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_right := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1970_c21_1af7_iftrue := resize(to_unsigned(0, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1955_c3_9fc5 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1955_c3_9fc5;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_374c_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c21_a00d_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_374c_left := VAR_phase;
     VAR_BIN_OP_DIV_uxn_opcodes_h_l1970_c35_bf62_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_DIV_uxn_opcodes_h_l1970_c35_bf62_right := t8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c21_a00d_left := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1961_l1953_l1958_l1972_DUPLICATE_21a0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1961_l1953_l1958_l1972_DUPLICATE_21a0_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1961_l1953_l1964_l1958_DUPLICATE_22d5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1961_l1953_l1964_l1958_DUPLICATE_22d5_return_output := result.u8_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1961_l1953_l1964_l1958_DUPLICATE_62fe LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1961_l1953_l1964_l1958_DUPLICATE_62fe_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1953_c6_f299] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_left;
     BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_return_output := BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1961_c11_a553] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_left;
     BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_return_output := BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1961_l1953_l1958_l1972_DUPLICATE_3e93 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1961_l1953_l1958_l1972_DUPLICATE_3e93_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1961_l1964_DUPLICATE_2fdb LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1961_l1964_DUPLICATE_2fdb_return_output := result.stack_address_sp_offset;

     -- BIN_OP_DIV[uxn_opcodes_h_l1970_c35_bf62] LATENCY=0
     -- Inputs
     BIN_OP_DIV_uxn_opcodes_h_l1970_c35_bf62_left <= VAR_BIN_OP_DIV_uxn_opcodes_h_l1970_c35_bf62_left;
     BIN_OP_DIV_uxn_opcodes_h_l1970_c35_bf62_right <= VAR_BIN_OP_DIV_uxn_opcodes_h_l1970_c35_bf62_right;
     -- Outputs
     VAR_BIN_OP_DIV_uxn_opcodes_h_l1970_c35_bf62_return_output := BIN_OP_DIV_uxn_opcodes_h_l1970_c35_bf62_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1972_c11_374c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1972_c11_374c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_374c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1972_c11_374c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_374c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_374c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1972_c11_374c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1958_c11_6068] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_left;
     BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_return_output := BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1961_l1964_l1958_l1972_DUPLICATE_3cd0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1961_l1964_l1958_l1972_DUPLICATE_3cd0_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1964_c11_3e14] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_left;
     BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_return_output := BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1970_c21_a00d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1970_c21_a00d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c21_a00d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1970_c21_a00d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c21_a00d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c21_a00d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1970_c21_a00d_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1967_c30_4d76] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_ins;
     sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_x;
     sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_return_output := sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_return_output;

     -- Submodule level 1
     VAR_MUX_uxn_opcodes_h_l1970_c21_1af7_iffalse := VAR_BIN_OP_DIV_uxn_opcodes_h_l1970_c35_bf62_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1953_c2_8dca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1953_c2_8dca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1953_c6_f299_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1958_c11_6068_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1961_c11_a553_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1964_c7_96da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1964_c11_3e14_return_output;
     VAR_MUX_uxn_opcodes_h_l1970_c21_1af7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c21_a00d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_374c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_374c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1972_c11_374c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1961_l1953_l1964_l1958_DUPLICATE_62fe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1961_l1953_l1964_l1958_DUPLICATE_62fe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1961_l1953_l1964_l1958_DUPLICATE_62fe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1961_l1953_l1964_l1958_DUPLICATE_62fe_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1961_l1964_l1958_l1972_DUPLICATE_3cd0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1961_l1964_l1958_l1972_DUPLICATE_3cd0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1961_l1964_l1958_l1972_DUPLICATE_3cd0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1961_l1964_l1958_l1972_DUPLICATE_3cd0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1961_l1953_l1958_l1972_DUPLICATE_21a0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1961_l1953_l1958_l1972_DUPLICATE_21a0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1961_l1953_l1958_l1972_DUPLICATE_21a0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1961_l1953_l1958_l1972_DUPLICATE_21a0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1961_l1953_l1958_l1972_DUPLICATE_3e93_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1961_l1953_l1958_l1972_DUPLICATE_3e93_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1961_l1953_l1958_l1972_DUPLICATE_3e93_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1961_l1953_l1958_l1972_DUPLICATE_3e93_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1961_l1964_DUPLICATE_2fdb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1961_l1964_DUPLICATE_2fdb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1961_l1953_l1964_l1958_DUPLICATE_22d5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1961_l1953_l1964_l1958_DUPLICATE_22d5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1961_l1953_l1964_l1958_DUPLICATE_22d5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1961_l1953_l1964_l1958_DUPLICATE_22d5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1967_c30_4d76_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1953_c1_fcb0] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1972_c7_9e83] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_return_output;

     -- n8_MUX[uxn_opcodes_h_l1964_c7_96da] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1964_c7_96da_cond <= VAR_n8_MUX_uxn_opcodes_h_l1964_c7_96da_cond;
     n8_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue;
     n8_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1964_c7_96da_return_output := n8_MUX_uxn_opcodes_h_l1964_c7_96da_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1972_c7_9e83] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1964_c7_96da] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1964_c7_96da] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1972_c7_9e83] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_return_output;

     -- t8_MUX[uxn_opcodes_h_l1961_c7_1b7a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond <= VAR_t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond;
     t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue;
     t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output := t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output;

     -- MUX[uxn_opcodes_h_l1970_c21_1af7] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1970_c21_1af7_cond <= VAR_MUX_uxn_opcodes_h_l1970_c21_1af7_cond;
     MUX_uxn_opcodes_h_l1970_c21_1af7_iftrue <= VAR_MUX_uxn_opcodes_h_l1970_c21_1af7_iftrue;
     MUX_uxn_opcodes_h_l1970_c21_1af7_iffalse <= VAR_MUX_uxn_opcodes_h_l1970_c21_1af7_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1970_c21_1af7_return_output := MUX_uxn_opcodes_h_l1970_c21_1af7_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue := VAR_MUX_uxn_opcodes_h_l1970_c21_1af7_return_output;
     VAR_printf_uxn_opcodes_h_l1954_c3_53b9_uxn_opcodes_h_l1954_c3_53b9_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1953_c1_fcb0_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1964_c7_96da_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1972_c7_9e83_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1972_c7_9e83_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1972_c7_9e83_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1964_c7_96da_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1964_c7_96da_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1964_c7_96da] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_return_output;

     -- t8_MUX[uxn_opcodes_h_l1958_c7_c9d8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond <= VAR_t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond;
     t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue;
     t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output := t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1964_c7_96da] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1961_c7_1b7a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1964_c7_96da] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1964_c7_96da] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_return_output := result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_return_output;

     -- printf_uxn_opcodes_h_l1954_c3_53b9[uxn_opcodes_h_l1954_c3_53b9] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1954_c3_53b9_uxn_opcodes_h_l1954_c3_53b9_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1954_c3_53b9_uxn_opcodes_h_l1954_c3_53b9_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1961_c7_1b7a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output;

     -- n8_MUX[uxn_opcodes_h_l1961_c7_1b7a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond <= VAR_n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond;
     n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue;
     n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output := n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1964_c7_96da_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1964_c7_96da_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1964_c7_96da_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1964_c7_96da_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1958_c7_c9d8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1961_c7_1b7a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1961_c7_1b7a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1961_c7_1b7a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output;

     -- n8_MUX[uxn_opcodes_h_l1958_c7_c9d8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond <= VAR_n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond;
     n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue;
     n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output := n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output;

     -- t8_MUX[uxn_opcodes_h_l1953_c2_8dca] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1953_c2_8dca_cond <= VAR_t8_MUX_uxn_opcodes_h_l1953_c2_8dca_cond;
     t8_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue;
     t8_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output := t8_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1961_c7_1b7a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output := result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1958_c7_c9d8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1961_c7_1b7a_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1958_c7_c9d8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output := result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1958_c7_c9d8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1953_c2_8dca] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1958_c7_c9d8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1958_c7_c9d8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1953_c2_8dca] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output;

     -- n8_MUX[uxn_opcodes_h_l1953_c2_8dca] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1953_c2_8dca_cond <= VAR_n8_MUX_uxn_opcodes_h_l1953_c2_8dca_cond;
     n8_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue;
     n8_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output := n8_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1958_c7_c9d8_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1953_c2_8dca] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1953_c2_8dca] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1953_c2_8dca] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output := result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1953_c2_8dca] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1978_l1949_DUPLICATE_1c81 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1978_l1949_DUPLICATE_1c81_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1953_c2_8dca_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1978_l1949_DUPLICATE_1c81_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1978_l1949_DUPLICATE_1c81_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
