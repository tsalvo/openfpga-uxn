-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 41
entity lit2_0CLK_4351dde2 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end lit2_0CLK_4351dde2;
architecture arch of lit2_0CLK_4351dde2 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal tmp8_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_tmp8_high : unsigned(7 downto 0);
signal REG_COMB_tmp8_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l219_c6_d2f3]
signal BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l219_c2_8e25]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l219_c2_8e25]
signal result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l219_c2_8e25]
signal result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l219_c2_8e25]
signal result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l219_c2_8e25]
signal result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l219_c2_8e25]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l219_c2_8e25]
signal result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l219_c2_8e25]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l219_c2_8e25]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l219_c2_8e25]
signal result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(0 downto 0);

-- tmp8_high_MUX[uxn_opcodes_h_l219_c2_8e25]
signal tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_cond : unsigned(0 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(7 downto 0);

-- tmp8_low_MUX[uxn_opcodes_h_l219_c2_8e25]
signal tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_cond : unsigned(0 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l232_c11_8a40]
signal BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l232_c7_2267]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l232_c7_2267]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l232_c7_2267]
signal result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l232_c7_2267]
signal result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l232_c7_2267]
signal result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l232_c7_2267]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l232_c7_2267]
signal result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_return_output : unsigned(0 downto 0);

-- tmp8_high_MUX[uxn_opcodes_h_l232_c7_2267]
signal tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_cond : unsigned(0 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_iftrue : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_iffalse : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_return_output : unsigned(7 downto 0);

-- tmp8_low_MUX[uxn_opcodes_h_l232_c7_2267]
signal tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_cond : unsigned(0 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_iftrue : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_iffalse : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_return_output : unsigned(7 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l234_c22_dc6a]
signal BIN_OP_PLUS_uxn_opcodes_h_l234_c22_dc6a_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l234_c22_dc6a_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l234_c22_dc6a_return_output : unsigned(16 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l236_c11_f7ea]
signal BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l236_c7_2fee]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l236_c7_2fee]
signal result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l236_c7_2fee]
signal result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l236_c7_2fee]
signal result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l236_c7_2fee]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l236_c7_2fee]
signal result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_return_output : unsigned(0 downto 0);

-- tmp8_high_MUX[uxn_opcodes_h_l236_c7_2fee]
signal tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_cond : unsigned(0 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_return_output : unsigned(7 downto 0);

-- tmp8_low_MUX[uxn_opcodes_h_l236_c7_2fee]
signal tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_cond : unsigned(0 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_return_output : unsigned(7 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l240_c22_307f]
signal BIN_OP_PLUS_uxn_opcodes_h_l240_c22_307f_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l240_c22_307f_right : unsigned(1 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l240_c22_307f_return_output : unsigned(16 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l244_c11_0743]
signal BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l244_c7_8db8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l244_c7_8db8]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l244_c7_8db8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l244_c7_8db8]
signal result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_return_output : unsigned(7 downto 0);

-- tmp8_low_MUX[uxn_opcodes_h_l244_c7_8db8]
signal tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_cond : unsigned(0 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_500b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_pc_updated := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.u16_value := ref_toks_4;
      base.is_ram_write := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_stack_write := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_stack_index_flipped := ref_toks_9;
      base.is_opc_done := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3
BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_left,
BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_right,
BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25
result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25
result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25
result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_cond,
result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25
result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_cond,
result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25
result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25
result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25
result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25
result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_return_output);

-- tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25
tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_cond,
tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue,
tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse,
tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_return_output);

-- tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25
tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_cond,
tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue,
tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse,
tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40
BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_left,
BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_right,
BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267
result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267
result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267
result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267
result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_cond,
result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267
result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_cond,
result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267
result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_return_output);

-- tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267
tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_cond,
tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_iftrue,
tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_iffalse,
tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_return_output);

-- tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267
tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_cond,
tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_iftrue,
tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_iffalse,
tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l234_c22_dc6a
BIN_OP_PLUS_uxn_opcodes_h_l234_c22_dc6a : entity work.BIN_OP_PLUS_uint16_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l234_c22_dc6a_left,
BIN_OP_PLUS_uxn_opcodes_h_l234_c22_dc6a_right,
BIN_OP_PLUS_uxn_opcodes_h_l234_c22_dc6a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea
BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_left,
BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_right,
BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee
result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee
result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee
result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_cond,
result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee
result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_cond,
result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee
result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_return_output);

-- tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee
tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_cond,
tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue,
tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse,
tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_return_output);

-- tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee
tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_cond,
tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue,
tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse,
tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l240_c22_307f
BIN_OP_PLUS_uxn_opcodes_h_l240_c22_307f : entity work.BIN_OP_PLUS_uint16_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l240_c22_307f_left,
BIN_OP_PLUS_uxn_opcodes_h_l240_c22_307f_right,
BIN_OP_PLUS_uxn_opcodes_h_l240_c22_307f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743
BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743_left,
BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743_right,
BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8
result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8
result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8
result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_cond,
result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_return_output);

-- tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8
tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_cond,
tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue,
tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse,
tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 previous_ram_read,
 -- Registers
 tmp8_high,
 tmp8_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_return_output,
 tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_return_output,
 tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_return_output,
 tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_return_output,
 tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l234_c22_dc6a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_return_output,
 tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_return_output,
 tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l240_c22_307f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_return_output,
 tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l228_c3_ffa2 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_cond : unsigned(0 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_cond : unsigned(0 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l233_c3_e674 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l232_c7_2267_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l234_c3_3e32 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_cond : unsigned(0 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_cond : unsigned(0 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l234_c22_dc6a_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l234_c22_dc6a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l234_c22_dc6a_return_output : unsigned(16 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l240_c3_469b : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_FALSE_INPUT_MUX_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l236_c7_2fee_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l241_c3_2893 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_cond : unsigned(0 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_cond : unsigned(0 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l240_c22_307f_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l240_c22_307f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l240_c22_307f_return_output : unsigned(16 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l247_c3_6627 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_cond : unsigned(0 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l232_l219_l244_DUPLICATE_7f6b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l232_l219_l244_DUPLICATE_80b4_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l232_l244_DUPLICATE_1b13_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l232_l236_DUPLICATE_4f30_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l232_l236_l244_DUPLICATE_72a2_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_500b_uxn_opcodes_h_l252_l214_DUPLICATE_76a8_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_tmp8_high : unsigned(7 downto 0);
variable REG_VAR_tmp8_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_tmp8_high := tmp8_high;
  REG_VAR_tmp8_low := tmp8_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_right := to_unsigned(2, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l228_c3_ffa2 := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l228_c3_ffa2;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l241_c3_2893 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l241_c3_2893;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743_right := to_unsigned(3, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l247_c3_6627 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l247_c3_6627;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l240_c22_307f_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_right := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l233_c3_e674 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l233_c3_e674;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l234_c22_dc6a_right := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l234_c22_dc6a_left := VAR_pc;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l240_c22_307f_left := VAR_pc;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue := VAR_previous_ram_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue := VAR_previous_ram_read;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue := VAR_previous_ram_read;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue := VAR_previous_ram_read;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue := tmp8_high;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_iftrue := tmp8_high;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse := tmp8_high;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue := tmp8_low;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_iftrue := tmp8_low;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue := tmp8_low;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse := tmp8_low;
     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l219_c2_8e25] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l219_c2_8e25_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l232_l236_l244_DUPLICATE_72a2 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l232_l236_l244_DUPLICATE_72a2_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l232_l244_DUPLICATE_1b13 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l232_l244_DUPLICATE_1b13_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l219_c6_d2f3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_left;
     BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_return_output := BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l232_l219_l244_DUPLICATE_80b4 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l232_l219_l244_DUPLICATE_80b4_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l232_l219_l244_DUPLICATE_7f6b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l232_l219_l244_DUPLICATE_7f6b_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l236_c11_f7ea] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_left;
     BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_return_output := BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l219_c2_8e25] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l219_c2_8e25_return_output := result.is_vram_write;

     -- result_u16_value_FALSE_INPUT_MUX_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d[uxn_opcodes_h_l236_c7_2fee] LATENCY=0
     VAR_result_u16_value_FALSE_INPUT_MUX_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l236_c7_2fee_return_output := result.u16_value;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l219_c2_8e25] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l219_c2_8e25_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l232_c11_8a40] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_left;
     BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_return_output := BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l232_l236_DUPLICATE_4f30 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l232_l236_DUPLICATE_4f30_return_output := result.is_stack_write;

     -- BIN_OP_PLUS[uxn_opcodes_h_l240_c22_307f] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l240_c22_307f_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l240_c22_307f_left;
     BIN_OP_PLUS_uxn_opcodes_h_l240_c22_307f_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l240_c22_307f_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l240_c22_307f_return_output := BIN_OP_PLUS_uxn_opcodes_h_l240_c22_307f_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l234_c22_dc6a] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l234_c22_dc6a_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l234_c22_dc6a_left;
     BIN_OP_PLUS_uxn_opcodes_h_l234_c22_dc6a_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l234_c22_dc6a_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l234_c22_dc6a_return_output := BIN_OP_PLUS_uxn_opcodes_h_l234_c22_dc6a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l244_c11_0743] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743_left;
     BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743_return_output := BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743_return_output;

     -- result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d[uxn_opcodes_h_l232_c7_2267] LATENCY=0
     VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l232_c7_2267_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_d2f3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_8a40_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_f7ea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_0743_return_output;
     VAR_result_u16_value_uxn_opcodes_h_l234_c3_3e32 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l234_c22_dc6a_return_output, 16);
     VAR_result_u16_value_uxn_opcodes_h_l240_c3_469b := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l240_c22_307f_return_output, 16);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l232_l236_l244_DUPLICATE_72a2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l232_l236_l244_DUPLICATE_72a2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l232_l236_l244_DUPLICATE_72a2_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l232_l244_DUPLICATE_1b13_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l232_l244_DUPLICATE_1b13_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l232_l236_DUPLICATE_4f30_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l232_l236_DUPLICATE_4f30_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l232_l219_l244_DUPLICATE_80b4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l232_l219_l244_DUPLICATE_80b4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l232_l219_l244_DUPLICATE_80b4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l232_l219_l244_DUPLICATE_7f6b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l232_l219_l244_DUPLICATE_7f6b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l232_l219_l244_DUPLICATE_7f6b_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l219_c2_8e25_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l219_c2_8e25_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l219_c2_8e25_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_iffalse := VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l232_c7_2267_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse := VAR_result_u16_value_FALSE_INPUT_MUX_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l236_c7_2fee_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_iftrue := VAR_result_u16_value_uxn_opcodes_h_l234_c3_3e32;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue := VAR_result_u16_value_uxn_opcodes_h_l240_c3_469b;
     -- result_is_vram_write_MUX[uxn_opcodes_h_l219_c2_8e25] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l244_c7_8db8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l236_c7_2fee] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_cond;
     result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_return_output := result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_return_output;

     -- tmp8_low_MUX[uxn_opcodes_h_l244_c7_8db8] LATENCY=0
     -- Inputs
     tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_cond <= VAR_tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_cond;
     tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue <= VAR_tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue;
     tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse <= VAR_tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse;
     -- Outputs
     VAR_tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_return_output := tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l236_c7_2fee] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l232_c7_2267] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l219_c2_8e25] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l219_c2_8e25] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l244_c7_8db8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l244_c7_8db8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_return_output := result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l244_c7_8db8] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_return_output;

     -- tmp8_high_MUX[uxn_opcodes_h_l236_c7_2fee] LATENCY=0
     -- Inputs
     tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_cond <= VAR_tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_cond;
     tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue <= VAR_tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue;
     tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse <= VAR_tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse;
     -- Outputs
     VAR_tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_return_output := tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_8db8_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_8db8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_2fee_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_2267_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_8db8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l236_c7_2fee_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l244_c7_8db8_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_iffalse := VAR_tmp8_high_MUX_uxn_opcodes_h_l236_c7_2fee_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse := VAR_tmp8_low_MUX_uxn_opcodes_h_l244_c7_8db8_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l236_c7_2fee] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_return_output;

     -- tmp8_low_MUX[uxn_opcodes_h_l236_c7_2fee] LATENCY=0
     -- Inputs
     tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_cond <= VAR_tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_cond;
     tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue <= VAR_tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue;
     tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse <= VAR_tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse;
     -- Outputs
     VAR_tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_return_output := tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l236_c7_2fee] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l236_c7_2fee] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l232_c7_2267] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_cond;
     result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_return_output := result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_return_output;

     -- tmp8_high_MUX[uxn_opcodes_h_l232_c7_2267] LATENCY=0
     -- Inputs
     tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_cond <= VAR_tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_cond;
     tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_iftrue <= VAR_tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_iftrue;
     tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_iffalse <= VAR_tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_iffalse;
     -- Outputs
     VAR_tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_return_output := tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l232_c7_2267] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l236_c7_2fee] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_cond;
     result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_return_output := result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l219_c2_8e25] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_2fee_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_2fee_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_2267_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_2fee_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l232_c7_2267_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l236_c7_2fee_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse := VAR_tmp8_high_MUX_uxn_opcodes_h_l232_c7_2267_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_iffalse := VAR_tmp8_low_MUX_uxn_opcodes_h_l236_c7_2fee_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l219_c2_8e25] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_return_output;

     -- tmp8_low_MUX[uxn_opcodes_h_l232_c7_2267] LATENCY=0
     -- Inputs
     tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_cond <= VAR_tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_cond;
     tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_iftrue <= VAR_tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_iftrue;
     tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_iffalse <= VAR_tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_iffalse;
     -- Outputs
     VAR_tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_return_output := tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_return_output;

     -- tmp8_high_MUX[uxn_opcodes_h_l219_c2_8e25] LATENCY=0
     -- Inputs
     tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_cond <= VAR_tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_cond;
     tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue <= VAR_tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue;
     tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse <= VAR_tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse;
     -- Outputs
     VAR_tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_return_output := tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l232_c7_2267] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_cond;
     result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_return_output := result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l219_c2_8e25] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_cond;
     result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_return_output := result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l232_c7_2267] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l232_c7_2267] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l232_c7_2267] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_2267_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_2267_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_2267_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l232_c7_2267_return_output;
     REG_VAR_tmp8_high := VAR_tmp8_high_MUX_uxn_opcodes_h_l219_c2_8e25_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse := VAR_tmp8_low_MUX_uxn_opcodes_h_l232_c7_2267_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l219_c2_8e25] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_cond;
     result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_return_output := result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l219_c2_8e25] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_return_output;

     -- tmp8_low_MUX[uxn_opcodes_h_l219_c2_8e25] LATENCY=0
     -- Inputs
     tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_cond <= VAR_tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_cond;
     tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue <= VAR_tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue;
     tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse <= VAR_tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse;
     -- Outputs
     VAR_tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_return_output := tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l219_c2_8e25] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l219_c2_8e25] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_return_output;

     -- Submodule level 5
     REG_VAR_tmp8_low := VAR_tmp8_low_MUX_uxn_opcodes_h_l219_c2_8e25_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_500b_uxn_opcodes_h_l252_l214_DUPLICATE_76a8 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_500b_uxn_opcodes_h_l252_l214_DUPLICATE_76a8_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_500b(
     result,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_8e25_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_8e25_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l219_c2_8e25_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l219_c2_8e25_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_8e25_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_8e25_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_8e25_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_8e25_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_8e25_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_8e25_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_500b_uxn_opcodes_h_l252_l214_DUPLICATE_76a8_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_500b_uxn_opcodes_h_l252_l214_DUPLICATE_76a8_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_tmp8_high <= REG_VAR_tmp8_high;
REG_COMB_tmp8_low <= REG_VAR_tmp8_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     tmp8_high <= REG_COMB_tmp8_high;
     tmp8_low <= REG_COMB_tmp8_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
