-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 57
entity sub_0CLK_edc09f97 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sub_0CLK_edc09f97;
architecture arch of sub_0CLK_edc09f97 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2685_c6_67cc]
signal BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2685_c2_858c]
signal n8_MUX_uxn_opcodes_h_l2685_c2_858c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2685_c2_858c_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2685_c2_858c]
signal t8_MUX_uxn_opcodes_h_l2685_c2_858c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2685_c2_858c_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2685_c2_858c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2685_c2_858c]
signal result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2685_c2_858c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2685_c2_858c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2685_c2_858c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2685_c2_858c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2690_c11_a415]
signal BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2690_c7_a426]
signal n8_MUX_uxn_opcodes_h_l2690_c7_a426_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2690_c7_a426_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2690_c7_a426]
signal t8_MUX_uxn_opcodes_h_l2690_c7_a426_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2690_c7_a426_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2690_c7_a426]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2690_c7_a426]
signal result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2690_c7_a426]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2690_c7_a426]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2690_c7_a426]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2690_c7_a426]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2693_c11_d833]
signal BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2693_c7_6858]
signal n8_MUX_uxn_opcodes_h_l2693_c7_6858_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2693_c7_6858_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2693_c7_6858]
signal t8_MUX_uxn_opcodes_h_l2693_c7_6858_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2693_c7_6858_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2693_c7_6858]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2693_c7_6858]
signal result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2693_c7_6858]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2693_c7_6858]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2693_c7_6858]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2693_c7_6858]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2697_c11_a8da]
signal BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2697_c7_9759]
signal n8_MUX_uxn_opcodes_h_l2697_c7_9759_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2697_c7_9759_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2697_c7_9759]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2697_c7_9759]
signal result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2697_c7_9759]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2697_c7_9759]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2697_c7_9759]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2697_c7_9759]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2700_c11_543b]
signal BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2700_c7_56c9]
signal n8_MUX_uxn_opcodes_h_l2700_c7_56c9_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2700_c7_56c9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2700_c7_56c9]
signal result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2700_c7_56c9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2700_c7_56c9]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2700_c7_56c9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2700_c7_56c9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l2703_c32_f8ef]
signal BIN_OP_AND_uxn_opcodes_h_l2703_c32_f8ef_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2703_c32_f8ef_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2703_c32_f8ef_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l2703_c32_5fe3]
signal BIN_OP_GT_uxn_opcodes_h_l2703_c32_5fe3_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l2703_c32_5fe3_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l2703_c32_5fe3_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l2703_c32_cf16]
signal MUX_uxn_opcodes_h_l2703_c32_cf16_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l2703_c32_cf16_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l2703_c32_cf16_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l2703_c32_cf16_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2705_c11_8bdf]
signal BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2705_c7_1b00]
signal result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2705_c7_1b00]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2705_c7_1b00]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2705_c7_1b00]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2705_c7_1b00]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output : unsigned(0 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_h_l2709_c24_e722]
signal BIN_OP_MINUS_uxn_opcodes_h_l2709_c24_e722_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2709_c24_e722_right : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2709_c24_e722_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2711_c11_2030]
signal BIN_OP_EQ_uxn_opcodes_h_l2711_c11_2030_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2711_c11_2030_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2711_c11_2030_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2711_c7_a376]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2711_c7_a376]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_value := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_sp_shift := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.is_opc_done := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc
BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_left,
BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_right,
BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_return_output);

-- n8_MUX_uxn_opcodes_h_l2685_c2_858c
n8_MUX_uxn_opcodes_h_l2685_c2_858c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2685_c2_858c_cond,
n8_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue,
n8_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse,
n8_MUX_uxn_opcodes_h_l2685_c2_858c_return_output);

-- t8_MUX_uxn_opcodes_h_l2685_c2_858c
t8_MUX_uxn_opcodes_h_l2685_c2_858c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2685_c2_858c_cond,
t8_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue,
t8_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse,
t8_MUX_uxn_opcodes_h_l2685_c2_858c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c
result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_cond,
result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c
result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c
result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c
result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415
BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_left,
BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_right,
BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_return_output);

-- n8_MUX_uxn_opcodes_h_l2690_c7_a426
n8_MUX_uxn_opcodes_h_l2690_c7_a426 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2690_c7_a426_cond,
n8_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue,
n8_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse,
n8_MUX_uxn_opcodes_h_l2690_c7_a426_return_output);

-- t8_MUX_uxn_opcodes_h_l2690_c7_a426
t8_MUX_uxn_opcodes_h_l2690_c7_a426 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2690_c7_a426_cond,
t8_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue,
t8_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse,
t8_MUX_uxn_opcodes_h_l2690_c7_a426_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426
result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426
result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_cond,
result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426
result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426
result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426
result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833
BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_left,
BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_right,
BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_return_output);

-- n8_MUX_uxn_opcodes_h_l2693_c7_6858
n8_MUX_uxn_opcodes_h_l2693_c7_6858 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2693_c7_6858_cond,
n8_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue,
n8_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse,
n8_MUX_uxn_opcodes_h_l2693_c7_6858_return_output);

-- t8_MUX_uxn_opcodes_h_l2693_c7_6858
t8_MUX_uxn_opcodes_h_l2693_c7_6858 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2693_c7_6858_cond,
t8_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue,
t8_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse,
t8_MUX_uxn_opcodes_h_l2693_c7_6858_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858
result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858
result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_cond,
result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858
result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858
result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858
result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da
BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_left,
BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_right,
BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_return_output);

-- n8_MUX_uxn_opcodes_h_l2697_c7_9759
n8_MUX_uxn_opcodes_h_l2697_c7_9759 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2697_c7_9759_cond,
n8_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue,
n8_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse,
n8_MUX_uxn_opcodes_h_l2697_c7_9759_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759
result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759
result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_cond,
result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759
result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759
result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759
result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b
BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_left,
BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_right,
BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_return_output);

-- n8_MUX_uxn_opcodes_h_l2700_c7_56c9
n8_MUX_uxn_opcodes_h_l2700_c7_56c9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2700_c7_56c9_cond,
n8_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue,
n8_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse,
n8_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9
result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9
result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_cond,
result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9
result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9
result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9
result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l2703_c32_f8ef
BIN_OP_AND_uxn_opcodes_h_l2703_c32_f8ef : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l2703_c32_f8ef_left,
BIN_OP_AND_uxn_opcodes_h_l2703_c32_f8ef_right,
BIN_OP_AND_uxn_opcodes_h_l2703_c32_f8ef_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l2703_c32_5fe3
BIN_OP_GT_uxn_opcodes_h_l2703_c32_5fe3 : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l2703_c32_5fe3_left,
BIN_OP_GT_uxn_opcodes_h_l2703_c32_5fe3_right,
BIN_OP_GT_uxn_opcodes_h_l2703_c32_5fe3_return_output);

-- MUX_uxn_opcodes_h_l2703_c32_cf16
MUX_uxn_opcodes_h_l2703_c32_cf16 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l2703_c32_cf16_cond,
MUX_uxn_opcodes_h_l2703_c32_cf16_iftrue,
MUX_uxn_opcodes_h_l2703_c32_cf16_iffalse,
MUX_uxn_opcodes_h_l2703_c32_cf16_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf
BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf_left,
BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf_right,
BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00
result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_cond,
result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00
result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00
result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00
result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l2709_c24_e722
BIN_OP_MINUS_uxn_opcodes_h_l2709_c24_e722 : entity work.BIN_OP_MINUS_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l2709_c24_e722_left,
BIN_OP_MINUS_uxn_opcodes_h_l2709_c24_e722_right,
BIN_OP_MINUS_uxn_opcodes_h_l2709_c24_e722_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2711_c11_2030
BIN_OP_EQ_uxn_opcodes_h_l2711_c11_2030 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2711_c11_2030_left,
BIN_OP_EQ_uxn_opcodes_h_l2711_c11_2030_right,
BIN_OP_EQ_uxn_opcodes_h_l2711_c11_2030_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376
result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376
result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_return_output,
 n8_MUX_uxn_opcodes_h_l2685_c2_858c_return_output,
 t8_MUX_uxn_opcodes_h_l2685_c2_858c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_return_output,
 n8_MUX_uxn_opcodes_h_l2690_c7_a426_return_output,
 t8_MUX_uxn_opcodes_h_l2690_c7_a426_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_return_output,
 n8_MUX_uxn_opcodes_h_l2693_c7_6858_return_output,
 t8_MUX_uxn_opcodes_h_l2693_c7_6858_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_return_output,
 n8_MUX_uxn_opcodes_h_l2697_c7_9759_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_return_output,
 n8_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output,
 BIN_OP_AND_uxn_opcodes_h_l2703_c32_f8ef_return_output,
 BIN_OP_GT_uxn_opcodes_h_l2703_c32_5fe3_return_output,
 MUX_uxn_opcodes_h_l2703_c32_cf16_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l2709_c24_e722_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2711_c11_2030_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2690_c7_a426_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2685_c2_858c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2685_c2_858c_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2690_c7_a426_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2685_c2_858c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2685_c2_858c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2687_c3_d7ac : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2693_c7_6858_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2690_c7_a426_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2693_c7_6858_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2690_c7_a426_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2691_c3_c478 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2697_c7_9759_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2693_c7_6858_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2693_c7_6858_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2695_c3_81b5 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2697_c7_9759_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2698_c3_1fab : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2700_c7_56c9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2703_c32_cf16_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2703_c32_cf16_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2703_c32_cf16_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2703_c32_f8ef_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2703_c32_f8ef_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2703_c32_f8ef_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2703_c32_5fe3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2703_c32_5fe3_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2703_c32_5fe3_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2703_c32_cf16_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2708_c3_f23f : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2709_c24_e722_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2709_c24_e722_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2709_c24_e722_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c11_2030_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c11_2030_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c11_2030_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_DUPLICATE_b147_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_l2705_DUPLICATE_6026_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2697_l2693_l2690_l2685_l2705_DUPLICATE_1971_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_l2711_DUPLICATE_e9b3_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2711_l2705_DUPLICATE_70b5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2700_l2705_DUPLICATE_4d1d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l2681_l2716_DUPLICATE_96cf_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2708_c3_f23f := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2708_c3_f23f;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2687_c3_d7ac := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2687_c3_d7ac;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2691_c3_c478 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2691_c3_c478;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l2703_c32_cf16_iffalse := resize(to_signed(-1, 2), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf_right := to_unsigned(5, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_AND_uxn_opcodes_h_l2703_c32_f8ef_right := to_unsigned(128, 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l2703_c32_cf16_iftrue := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_BIN_OP_GT_uxn_opcodes_h_l2703_c32_5fe3_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c11_2030_right := to_unsigned(6, 3);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2695_c3_81b5 := resize(to_unsigned(2, 2), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2695_c3_81b5;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2698_c3_1fab := resize(to_unsigned(2, 2), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2698_c3_1fab;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_BIN_OP_AND_uxn_opcodes_h_l2703_c32_f8ef_left := VAR_ins;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2709_c24_e722_left := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c11_2030_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2709_c24_e722_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2705_c11_8bdf] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf_left;
     BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf_return_output := BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf_return_output;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_DUPLICATE_b147 LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_DUPLICATE_b147_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_l2711_DUPLICATE_e9b3 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_l2711_DUPLICATE_e9b3_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2700_l2705_DUPLICATE_4d1d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2700_l2705_DUPLICATE_4d1d_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2700_c11_543b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_left;
     BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_return_output := BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l2703_c32_f8ef] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l2703_c32_f8ef_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l2703_c32_f8ef_left;
     BIN_OP_AND_uxn_opcodes_h_l2703_c32_f8ef_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l2703_c32_f8ef_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l2703_c32_f8ef_return_output := BIN_OP_AND_uxn_opcodes_h_l2703_c32_f8ef_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2685_c6_67cc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_left;
     BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_return_output := BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_l2705_DUPLICATE_6026 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_l2705_DUPLICATE_6026_return_output := result.stack_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2697_c11_a8da] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_left;
     BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_return_output := BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2693_c11_d833] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_left;
     BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_return_output := BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_return_output;

     -- BIN_OP_MINUS[uxn_opcodes_h_l2709_c24_e722] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l2709_c24_e722_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2709_c24_e722_left;
     BIN_OP_MINUS_uxn_opcodes_h_l2709_c24_e722_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2709_c24_e722_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2709_c24_e722_return_output := BIN_OP_MINUS_uxn_opcodes_h_l2709_c24_e722_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2690_c11_a415] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_left;
     BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_return_output := BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2711_l2705_DUPLICATE_70b5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2711_l2705_DUPLICATE_70b5_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2697_l2693_l2690_l2685_l2705_DUPLICATE_1971 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2697_l2693_l2690_l2685_l2705_DUPLICATE_1971_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2711_c11_2030] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2711_c11_2030_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c11_2030_left;
     BIN_OP_EQ_uxn_opcodes_h_l2711_c11_2030_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c11_2030_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c11_2030_return_output := BIN_OP_EQ_uxn_opcodes_h_l2711_c11_2030_return_output;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l2703_c32_5fe3_left := VAR_BIN_OP_AND_uxn_opcodes_h_l2703_c32_f8ef_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2685_c2_858c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2685_c2_858c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2685_c6_67cc_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2690_c7_a426_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2690_c7_a426_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2690_c11_a415_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2693_c7_6858_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2693_c7_6858_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2693_c11_d833_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2697_c7_9759_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2697_c11_a8da_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2700_c7_56c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2700_c11_543b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2705_c11_8bdf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c11_2030_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2711_c11_2030_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue := VAR_BIN_OP_MINUS_uxn_opcodes_h_l2709_c24_e722_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_DUPLICATE_b147_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_DUPLICATE_b147_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_DUPLICATE_b147_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_DUPLICATE_b147_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_DUPLICATE_b147_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2711_l2705_DUPLICATE_70b5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2711_l2705_DUPLICATE_70b5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2711_l2705_DUPLICATE_70b5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2711_l2705_DUPLICATE_70b5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2711_l2705_DUPLICATE_70b5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2711_l2705_DUPLICATE_70b5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2697_l2693_l2690_l2685_l2705_DUPLICATE_1971_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2697_l2693_l2690_l2685_l2705_DUPLICATE_1971_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2697_l2693_l2690_l2685_l2705_DUPLICATE_1971_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2697_l2693_l2690_l2685_l2705_DUPLICATE_1971_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2697_l2693_l2690_l2685_l2705_DUPLICATE_1971_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_l2711_DUPLICATE_e9b3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_l2711_DUPLICATE_e9b3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_l2711_DUPLICATE_e9b3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_l2711_DUPLICATE_e9b3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_l2711_DUPLICATE_e9b3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_l2711_DUPLICATE_e9b3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2700_l2705_DUPLICATE_4d1d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2700_l2705_DUPLICATE_4d1d_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_l2705_DUPLICATE_6026_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_l2705_DUPLICATE_6026_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_l2705_DUPLICATE_6026_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_l2705_DUPLICATE_6026_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_l2705_DUPLICATE_6026_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2700_l2697_l2693_l2690_l2685_l2705_DUPLICATE_6026_return_output;
     -- n8_MUX[uxn_opcodes_h_l2700_c7_56c9] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2700_c7_56c9_cond <= VAR_n8_MUX_uxn_opcodes_h_l2700_c7_56c9_cond;
     n8_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue;
     n8_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output := n8_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2705_c7_1b00] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output := result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2711_c7_a376] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_return_output;

     -- t8_MUX[uxn_opcodes_h_l2693_c7_6858] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2693_c7_6858_cond <= VAR_t8_MUX_uxn_opcodes_h_l2693_c7_6858_cond;
     t8_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue;
     t8_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2693_c7_6858_return_output := t8_MUX_uxn_opcodes_h_l2693_c7_6858_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2705_c7_1b00] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l2703_c32_5fe3] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l2703_c32_5fe3_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l2703_c32_5fe3_left;
     BIN_OP_GT_uxn_opcodes_h_l2703_c32_5fe3_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l2703_c32_5fe3_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l2703_c32_5fe3_return_output := BIN_OP_GT_uxn_opcodes_h_l2703_c32_5fe3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2705_c7_1b00] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2711_c7_a376] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l2703_c32_cf16_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l2703_c32_5fe3_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2711_c7_a376_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2711_c7_a376_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2693_c7_6858_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2700_c7_56c9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output;

     -- MUX[uxn_opcodes_h_l2703_c32_cf16] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l2703_c32_cf16_cond <= VAR_MUX_uxn_opcodes_h_l2703_c32_cf16_cond;
     MUX_uxn_opcodes_h_l2703_c32_cf16_iftrue <= VAR_MUX_uxn_opcodes_h_l2703_c32_cf16_iftrue;
     MUX_uxn_opcodes_h_l2703_c32_cf16_iffalse <= VAR_MUX_uxn_opcodes_h_l2703_c32_cf16_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l2703_c32_cf16_return_output := MUX_uxn_opcodes_h_l2703_c32_cf16_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2700_c7_56c9] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output := result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2705_c7_1b00] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2705_c7_1b00] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output;

     -- t8_MUX[uxn_opcodes_h_l2690_c7_a426] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2690_c7_a426_cond <= VAR_t8_MUX_uxn_opcodes_h_l2690_c7_a426_cond;
     t8_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue;
     t8_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2690_c7_a426_return_output := t8_MUX_uxn_opcodes_h_l2690_c7_a426_return_output;

     -- n8_MUX[uxn_opcodes_h_l2697_c7_9759] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2697_c7_9759_cond <= VAR_n8_MUX_uxn_opcodes_h_l2697_c7_9759_cond;
     n8_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue;
     n8_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2697_c7_9759_return_output := n8_MUX_uxn_opcodes_h_l2697_c7_9759_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2700_c7_56c9] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue := VAR_MUX_uxn_opcodes_h_l2703_c32_cf16_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2697_c7_9759_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2705_c7_1b00_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2690_c7_a426_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2700_c7_56c9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2700_c7_56c9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2697_c7_9759] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_return_output := result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2697_c7_9759] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2700_c7_56c9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2697_c7_9759] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_return_output;

     -- t8_MUX[uxn_opcodes_h_l2685_c2_858c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2685_c2_858c_cond <= VAR_t8_MUX_uxn_opcodes_h_l2685_c2_858c_cond;
     t8_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue;
     t8_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2685_c2_858c_return_output := t8_MUX_uxn_opcodes_h_l2685_c2_858c_return_output;

     -- n8_MUX[uxn_opcodes_h_l2693_c7_6858] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2693_c7_6858_cond <= VAR_n8_MUX_uxn_opcodes_h_l2693_c7_6858_cond;
     n8_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue;
     n8_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2693_c7_6858_return_output := n8_MUX_uxn_opcodes_h_l2693_c7_6858_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2693_c7_6858_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2697_c7_9759_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2700_c7_56c9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2697_c7_9759_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2697_c7_9759_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2685_c2_858c_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2693_c7_6858] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_return_output;

     -- n8_MUX[uxn_opcodes_h_l2690_c7_a426] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2690_c7_a426_cond <= VAR_n8_MUX_uxn_opcodes_h_l2690_c7_a426_cond;
     n8_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue;
     n8_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2690_c7_a426_return_output := n8_MUX_uxn_opcodes_h_l2690_c7_a426_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2697_c7_9759] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2697_c7_9759] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2697_c7_9759] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2693_c7_6858] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_return_output := result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2693_c7_6858] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2690_c7_a426_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2697_c7_9759_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2693_c7_6858_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2697_c7_9759_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2697_c7_9759_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2693_c7_6858_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2693_c7_6858_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2693_c7_6858] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_return_output;

     -- n8_MUX[uxn_opcodes_h_l2685_c2_858c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2685_c2_858c_cond <= VAR_n8_MUX_uxn_opcodes_h_l2685_c2_858c_cond;
     n8_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue;
     n8_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2685_c2_858c_return_output := n8_MUX_uxn_opcodes_h_l2685_c2_858c_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2690_c7_a426] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_return_output := result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2693_c7_6858] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2690_c7_a426] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2690_c7_a426] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2693_c7_6858] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2685_c2_858c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2693_c7_6858_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2690_c7_a426_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2693_c7_6858_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2693_c7_6858_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2690_c7_a426_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2690_c7_a426_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2690_c7_a426] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2685_c2_858c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2685_c2_858c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2690_c7_a426] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2690_c7_a426] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2685_c2_858c] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_return_output := result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_return_output;

     -- Submodule level 7
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2690_c7_a426_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2690_c7_a426_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2690_c7_a426_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2685_c2_858c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2685_c2_858c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2685_c2_858c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_return_output;

     -- Submodule level 8
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l2681_l2716_DUPLICATE_96cf LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l2681_l2716_DUPLICATE_96cf_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2685_c2_858c_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2685_c2_858c_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2685_c2_858c_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2685_c2_858c_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2685_c2_858c_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2685_c2_858c_return_output);

     -- Submodule level 9
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l2681_l2716_DUPLICATE_96cf_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l2681_l2716_DUPLICATE_96cf_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
