-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 37
entity dup_0CLK_6be78140 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dup_0CLK_6be78140;
architecture arch of dup_0CLK_6be78140 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2953_c6_6b7a]
signal BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2953_c1_267e]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2953_c2_c39e]
signal t8_MUX_uxn_opcodes_h_l2953_c2_c39e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2953_c2_c39e]
signal result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2953_c2_c39e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2953_c2_c39e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2953_c2_c39e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2953_c2_c39e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2953_c2_c39e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output : unsigned(3 downto 0);

-- printf_uxn_opcodes_h_l2954_c3_b3d9[uxn_opcodes_h_l2954_c3_b3d9]
signal printf_uxn_opcodes_h_l2954_c3_b3d9_uxn_opcodes_h_l2954_c3_b3d9_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2958_c11_331b]
signal BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2958_c7_e66b]
signal t8_MUX_uxn_opcodes_h_l2958_c7_e66b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2958_c7_e66b]
signal result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2958_c7_e66b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2958_c7_e66b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2958_c7_e66b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2958_c7_e66b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2958_c7_e66b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2961_c11_9be6]
signal BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2961_c7_ef0d]
signal t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2961_c7_ef0d]
signal result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2961_c7_ef0d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2961_c7_ef0d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2961_c7_ef0d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2961_c7_ef0d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2961_c7_ef0d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output : unsigned(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2964_c30_b989]
signal sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2969_c11_f940]
signal BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2969_c7_16a3]
signal result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2969_c7_16a3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2969_c7_16a3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2969_c7_16a3]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2969_c7_16a3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2974_c11_944c]
signal BIN_OP_EQ_uxn_opcodes_h_l2974_c11_944c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2974_c11_944c_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2974_c11_944c_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2974_c7_0251]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2974_c7_0251]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_25e8( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.is_sp_shift := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a
BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_left,
BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_right,
BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_return_output);

-- t8_MUX_uxn_opcodes_h_l2953_c2_c39e
t8_MUX_uxn_opcodes_h_l2953_c2_c39e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2953_c2_c39e_cond,
t8_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue,
t8_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse,
t8_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e
result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_cond,
result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e
result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e
result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e
result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e
result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output);

-- printf_uxn_opcodes_h_l2954_c3_b3d9_uxn_opcodes_h_l2954_c3_b3d9
printf_uxn_opcodes_h_l2954_c3_b3d9_uxn_opcodes_h_l2954_c3_b3d9 : entity work.printf_uxn_opcodes_h_l2954_c3_b3d9_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2954_c3_b3d9_uxn_opcodes_h_l2954_c3_b3d9_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b
BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_left,
BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_right,
BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_return_output);

-- t8_MUX_uxn_opcodes_h_l2958_c7_e66b
t8_MUX_uxn_opcodes_h_l2958_c7_e66b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2958_c7_e66b_cond,
t8_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue,
t8_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse,
t8_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b
result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_cond,
result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b
result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b
result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b
result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b
result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6
BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_left,
BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_right,
BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_return_output);

-- t8_MUX_uxn_opcodes_h_l2961_c7_ef0d
t8_MUX_uxn_opcodes_h_l2961_c7_ef0d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond,
t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue,
t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse,
t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d
result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond,
result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d
result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d
result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d
result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d
result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2964_c30_b989
sp_relative_shift_uxn_opcodes_h_l2964_c30_b989 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_ins,
sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_x,
sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_y,
sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940
BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940_left,
BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940_right,
BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3
result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_cond,
result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3
result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3
result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3
result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2974_c11_944c
BIN_OP_EQ_uxn_opcodes_h_l2974_c11_944c : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2974_c11_944c_left,
BIN_OP_EQ_uxn_opcodes_h_l2974_c11_944c_right,
BIN_OP_EQ_uxn_opcodes_h_l2974_c11_944c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251
result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251
result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_return_output,
 t8_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_return_output,
 t8_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_return_output,
 t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output,
 sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2974_c11_944c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2953_c2_c39e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2955_c3_da5a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2954_c3_b3d9_uxn_opcodes_h_l2954_c3_b3d9_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2958_c7_e66b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2959_c3_4334 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2966_c3_07d3 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2971_c3_6806 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2969_c7_16a3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2974_c11_944c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2974_c11_944c_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2974_c11_944c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2953_l2969_l2958_DUPLICATE_920b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2961_l2953_l2958_DUPLICATE_70ae_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2953_l2969_l2958_l2974_DUPLICATE_4e13_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2953_l2969_l2958_DUPLICATE_1200_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2961_l2969_l2958_l2974_DUPLICATE_86ce_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l2949_l2979_DUPLICATE_8072_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2974_c11_944c_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2959_c3_4334 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2959_c3_4334;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2966_c3_07d3 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2966_c3_07d3;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2955_c3_da5a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2955_c3_da5a;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2971_c3_6806 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2971_c3_6806;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2974_c11_944c_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse := t8;
     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2961_l2953_l2958_DUPLICATE_70ae LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2961_l2953_l2958_DUPLICATE_70ae_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2969_c11_f940] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940_left;
     BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940_return_output := BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2953_l2969_l2958_DUPLICATE_1200 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2953_l2969_l2958_DUPLICATE_1200_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2974_c11_944c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2974_c11_944c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2974_c11_944c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2974_c11_944c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2974_c11_944c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2974_c11_944c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2974_c11_944c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2953_c6_6b7a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2969_c7_16a3] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2969_c7_16a3_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2961_l2969_l2958_l2974_DUPLICATE_86ce LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2961_l2969_l2958_l2974_DUPLICATE_86ce_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2958_c11_331b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_left;
     BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_return_output := BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2953_l2969_l2958_l2974_DUPLICATE_4e13 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2953_l2969_l2958_l2974_DUPLICATE_4e13_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2953_l2969_l2958_DUPLICATE_920b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2953_l2969_l2958_DUPLICATE_920b_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2961_c11_9be6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_left;
     BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_return_output := BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2964_c30_b989] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_ins;
     sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_x;
     sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_return_output := sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2953_c2_c39e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2953_c6_6b7a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2958_c7_e66b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2958_c11_331b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2961_c11_9be6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2969_c11_f940_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2974_c11_944c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2974_c11_944c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2961_l2953_l2958_DUPLICATE_70ae_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2961_l2953_l2958_DUPLICATE_70ae_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2961_l2953_l2958_DUPLICATE_70ae_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2961_l2969_l2958_l2974_DUPLICATE_86ce_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2961_l2969_l2958_l2974_DUPLICATE_86ce_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2961_l2969_l2958_l2974_DUPLICATE_86ce_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2961_l2969_l2958_l2974_DUPLICATE_86ce_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2953_l2969_l2958_DUPLICATE_1200_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2953_l2969_l2958_DUPLICATE_1200_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2953_l2969_l2958_DUPLICATE_1200_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2953_l2969_l2958_l2974_DUPLICATE_4e13_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2953_l2969_l2958_l2974_DUPLICATE_4e13_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2953_l2969_l2958_l2974_DUPLICATE_4e13_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2953_l2969_l2958_l2974_DUPLICATE_4e13_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2953_l2969_l2958_DUPLICATE_920b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2953_l2969_l2958_DUPLICATE_920b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2953_l2969_l2958_DUPLICATE_920b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2969_c7_16a3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2964_c30_b989_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2974_c7_0251] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2969_c7_16a3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2974_c7_0251] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_return_output;

     -- t8_MUX[uxn_opcodes_h_l2961_c7_ef0d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond <= VAR_t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond;
     t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue;
     t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output := t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2969_c7_16a3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output := result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2969_c7_16a3] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2953_c1_267e] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2961_c7_ef0d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l2954_c3_b3d9_uxn_opcodes_h_l2954_c3_b3d9_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2953_c1_267e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2974_c7_0251_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2974_c7_0251_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2969_c7_16a3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output;

     -- printf_uxn_opcodes_h_l2954_c3_b3d9[uxn_opcodes_h_l2954_c3_b3d9] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2954_c3_b3d9_uxn_opcodes_h_l2954_c3_b3d9_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2954_c3_b3d9_uxn_opcodes_h_l2954_c3_b3d9_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2961_c7_ef0d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2969_c7_16a3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2961_c7_ef0d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output := result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2961_c7_ef0d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2958_c7_e66b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output;

     -- t8_MUX[uxn_opcodes_h_l2958_c7_e66b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2958_c7_e66b_cond <= VAR_t8_MUX_uxn_opcodes_h_l2958_c7_e66b_cond;
     t8_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue;
     t8_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output := t8_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2969_c7_16a3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2961_c7_ef0d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output;

     -- t8_MUX[uxn_opcodes_h_l2953_c2_c39e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2953_c2_c39e_cond <= VAR_t8_MUX_uxn_opcodes_h_l2953_c2_c39e_cond;
     t8_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue;
     t8_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output := t8_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2958_c7_e66b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2958_c7_e66b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output := result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2953_c2_c39e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2961_c7_ef0d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2958_c7_e66b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2961_c7_ef0d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2958_c7_e66b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2953_c2_c39e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2958_c7_e66b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2953_c2_c39e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output := result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2953_c2_c39e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2958_c7_e66b_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2953_c2_c39e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2953_c2_c39e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l2949_l2979_DUPLICATE_8072 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l2949_l2979_DUPLICATE_8072_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_25e8(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2953_c2_c39e_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l2949_l2979_DUPLICATE_8072_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l2949_l2979_DUPLICATE_8072_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
