-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity eor_0CLK_64d180f1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end eor_0CLK_64d180f1;
architecture arch of eor_0CLK_64d180f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1077_c6_07a2]
signal BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1077_c2_8c24]
signal n8_MUX_uxn_opcodes_h_l1077_c2_8c24_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1077_c2_8c24]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1077_c2_8c24]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1077_c2_8c24]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1077_c2_8c24]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1077_c2_8c24]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1077_c2_8c24]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1077_c2_8c24]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1077_c2_8c24]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1077_c2_8c24]
signal result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1077_c2_8c24]
signal t8_MUX_uxn_opcodes_h_l1077_c2_8c24_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1090_c11_6858]
signal BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1090_c7_3f35]
signal n8_MUX_uxn_opcodes_h_l1090_c7_3f35_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1090_c7_3f35]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1090_c7_3f35]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1090_c7_3f35]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1090_c7_3f35]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1090_c7_3f35]
signal result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1090_c7_3f35]
signal t8_MUX_uxn_opcodes_h_l1090_c7_3f35_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1093_c11_a1e8]
signal BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1093_c7_ca31]
signal n8_MUX_uxn_opcodes_h_l1093_c7_ca31_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1093_c7_ca31]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1093_c7_ca31]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1093_c7_ca31]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1093_c7_ca31]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1093_c7_ca31]
signal result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1093_c7_ca31]
signal t8_MUX_uxn_opcodes_h_l1093_c7_ca31_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1096_c11_af3d]
signal BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1096_c7_e9f8]
signal n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1096_c7_e9f8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1096_c7_e9f8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1096_c7_e9f8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1096_c7_e9f8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1096_c7_e9f8]
signal result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1098_c30_a1c1]
signal sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_return_output : signed(3 downto 0);

-- BIN_OP_XOR[uxn_opcodes_h_l1101_c21_e4ec]
signal BIN_OP_XOR_uxn_opcodes_h_l1101_c21_e4ec_left : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1101_c21_e4ec_right : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1101_c21_e4ec_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_04b4( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.is_stack_index_flipped := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.u8_value := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2
BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_left,
BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_right,
BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_return_output);

-- n8_MUX_uxn_opcodes_h_l1077_c2_8c24
n8_MUX_uxn_opcodes_h_l1077_c2_8c24 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1077_c2_8c24_cond,
n8_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue,
n8_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse,
n8_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24
result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24
result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24
result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24
result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24
result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24
result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24
result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_cond,
result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output);

-- t8_MUX_uxn_opcodes_h_l1077_c2_8c24
t8_MUX_uxn_opcodes_h_l1077_c2_8c24 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1077_c2_8c24_cond,
t8_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue,
t8_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse,
t8_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858
BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_left,
BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_right,
BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_return_output);

-- n8_MUX_uxn_opcodes_h_l1090_c7_3f35
n8_MUX_uxn_opcodes_h_l1090_c7_3f35 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1090_c7_3f35_cond,
n8_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue,
n8_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse,
n8_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35
result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35
result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35
result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35
result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_cond,
result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output);

-- t8_MUX_uxn_opcodes_h_l1090_c7_3f35
t8_MUX_uxn_opcodes_h_l1090_c7_3f35 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1090_c7_3f35_cond,
t8_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue,
t8_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse,
t8_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8
BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_left,
BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_right,
BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_return_output);

-- n8_MUX_uxn_opcodes_h_l1093_c7_ca31
n8_MUX_uxn_opcodes_h_l1093_c7_ca31 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1093_c7_ca31_cond,
n8_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue,
n8_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse,
n8_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31
result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31
result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31
result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31
result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_cond,
result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output);

-- t8_MUX_uxn_opcodes_h_l1093_c7_ca31
t8_MUX_uxn_opcodes_h_l1093_c7_ca31 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1093_c7_ca31_cond,
t8_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue,
t8_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse,
t8_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d
BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d_left,
BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d_right,
BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d_return_output);

-- n8_MUX_uxn_opcodes_h_l1096_c7_e9f8
n8_MUX_uxn_opcodes_h_l1096_c7_e9f8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond,
n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue,
n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse,
n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8
result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8
result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8
result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8
result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond,
result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1
sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_ins,
sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_x,
sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_y,
sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_return_output);

-- BIN_OP_XOR_uxn_opcodes_h_l1101_c21_e4ec
BIN_OP_XOR_uxn_opcodes_h_l1101_c21_e4ec : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_XOR_uxn_opcodes_h_l1101_c21_e4ec_left,
BIN_OP_XOR_uxn_opcodes_h_l1101_c21_e4ec_right,
BIN_OP_XOR_uxn_opcodes_h_l1101_c21_e4ec_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_return_output,
 n8_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output,
 t8_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_return_output,
 n8_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output,
 t8_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_return_output,
 n8_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output,
 t8_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d_return_output,
 n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output,
 sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_return_output,
 BIN_OP_XOR_uxn_opcodes_h_l1101_c21_e4ec_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1077_c2_8c24_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1077_c2_8c24_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1087_c3_1770 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1077_c2_8c24_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1082_c3_f04e : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1077_c2_8c24_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1077_c2_8c24_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1077_c2_8c24_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1090_c7_3f35_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1091_c3_bf85 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1090_c7_3f35_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1093_c7_ca31_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1093_c7_ca31_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1100_c3_1094 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1101_c21_e4ec_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1101_c21_e4ec_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1101_c21_e4ec_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1077_l1096_l1090_l1093_DUPLICATE_7b6e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1096_l1090_l1093_DUPLICATE_db24_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1096_l1090_l1093_DUPLICATE_2d5f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1096_l1090_l1093_DUPLICATE_36ea_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1096_l1093_DUPLICATE_ceda_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l1105_l1073_DUPLICATE_c0e4_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1082_c3_f04e := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1082_c3_f04e;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_y := resize(to_signed(-1, 2), 4);
     VAR_sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_right := to_unsigned(2, 2);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1087_c3_1770 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1087_c3_1770;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1100_c3_1094 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1100_c3_1094;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1091_c3_bf85 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1091_c3_bf85;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d_left := VAR_phase;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1101_c21_e4ec_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1101_c21_e4ec_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse := t8;
     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1077_c2_8c24] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1077_c2_8c24_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l1093_c11_a1e8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_left;
     BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_return_output := BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1077_c2_8c24] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1077_c2_8c24_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1077_l1096_l1090_l1093_DUPLICATE_7b6e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1077_l1096_l1090_l1093_DUPLICATE_7b6e_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1090_c11_6858] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_left;
     BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_return_output := BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1077_c2_8c24] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1077_c2_8c24_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1096_l1090_l1093_DUPLICATE_36ea LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1096_l1090_l1093_DUPLICATE_36ea_return_output := result.is_stack_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1077_c2_8c24] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1077_c2_8c24_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1096_l1093_DUPLICATE_ceda LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1096_l1093_DUPLICATE_ceda_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1077_c6_07a2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_left;
     BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_return_output := BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1096_l1090_l1093_DUPLICATE_db24 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1096_l1090_l1093_DUPLICATE_db24_return_output := result.sp_relative_shift;

     -- sp_relative_shift[uxn_opcodes_h_l1098_c30_a1c1] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_ins;
     sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_x;
     sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_return_output := sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_return_output;

     -- BIN_OP_XOR[uxn_opcodes_h_l1101_c21_e4ec] LATENCY=0
     -- Inputs
     BIN_OP_XOR_uxn_opcodes_h_l1101_c21_e4ec_left <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1101_c21_e4ec_left;
     BIN_OP_XOR_uxn_opcodes_h_l1101_c21_e4ec_right <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1101_c21_e4ec_right;
     -- Outputs
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1101_c21_e4ec_return_output := BIN_OP_XOR_uxn_opcodes_h_l1101_c21_e4ec_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1096_l1090_l1093_DUPLICATE_2d5f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1096_l1090_l1093_DUPLICATE_2d5f_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1096_c11_af3d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1077_c2_8c24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1077_c2_8c24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1077_c6_07a2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1090_c7_3f35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1090_c7_3f35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1090_c11_6858_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1093_c7_ca31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1093_c7_ca31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1093_c11_a1e8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1096_c11_af3d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue := VAR_BIN_OP_XOR_uxn_opcodes_h_l1101_c21_e4ec_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1096_l1090_l1093_DUPLICATE_db24_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1096_l1090_l1093_DUPLICATE_db24_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1096_l1090_l1093_DUPLICATE_db24_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1096_l1090_l1093_DUPLICATE_2d5f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1096_l1090_l1093_DUPLICATE_2d5f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1096_l1090_l1093_DUPLICATE_2d5f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1096_l1090_l1093_DUPLICATE_36ea_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1096_l1090_l1093_DUPLICATE_36ea_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1096_l1090_l1093_DUPLICATE_36ea_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1096_l1093_DUPLICATE_ceda_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1096_l1093_DUPLICATE_ceda_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1077_l1096_l1090_l1093_DUPLICATE_7b6e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1077_l1096_l1090_l1093_DUPLICATE_7b6e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1077_l1096_l1090_l1093_DUPLICATE_7b6e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1077_l1096_l1090_l1093_DUPLICATE_7b6e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1077_c2_8c24_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1077_c2_8c24_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1077_c2_8c24_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1077_c2_8c24_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1098_c30_a1c1_return_output;
     -- n8_MUX[uxn_opcodes_h_l1096_c7_e9f8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond <= VAR_n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond;
     n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue;
     n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output := n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1077_c2_8c24] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1096_c7_e9f8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1096_c7_e9f8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1077_c2_8c24] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1077_c2_8c24] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1096_c7_e9f8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1096_c7_e9f8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output := result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1077_c2_8c24] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output;

     -- t8_MUX[uxn_opcodes_h_l1093_c7_ca31] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1093_c7_ca31_cond <= VAR_t8_MUX_uxn_opcodes_h_l1093_c7_ca31_cond;
     t8_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue;
     t8_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output := t8_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1096_c7_e9f8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1096_c7_e9f8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1093_c7_ca31] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output := result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output;

     -- n8_MUX[uxn_opcodes_h_l1093_c7_ca31] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1093_c7_ca31_cond <= VAR_n8_MUX_uxn_opcodes_h_l1093_c7_ca31_cond;
     n8_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue;
     n8_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output := n8_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1093_c7_ca31] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1093_c7_ca31] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output;

     -- t8_MUX[uxn_opcodes_h_l1090_c7_3f35] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1090_c7_3f35_cond <= VAR_t8_MUX_uxn_opcodes_h_l1090_c7_3f35_cond;
     t8_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue;
     t8_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output := t8_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1093_c7_ca31] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1093_c7_ca31] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1093_c7_ca31_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1090_c7_3f35] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1090_c7_3f35] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1090_c7_3f35] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output;

     -- n8_MUX[uxn_opcodes_h_l1090_c7_3f35] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1090_c7_3f35_cond <= VAR_n8_MUX_uxn_opcodes_h_l1090_c7_3f35_cond;
     n8_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue;
     n8_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output := n8_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1090_c7_3f35] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1090_c7_3f35] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output := result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output;

     -- t8_MUX[uxn_opcodes_h_l1077_c2_8c24] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1077_c2_8c24_cond <= VAR_t8_MUX_uxn_opcodes_h_l1077_c2_8c24_cond;
     t8_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue;
     t8_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output := t8_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1090_c7_3f35_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output;
     -- n8_MUX[uxn_opcodes_h_l1077_c2_8c24] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1077_c2_8c24_cond <= VAR_n8_MUX_uxn_opcodes_h_l1077_c2_8c24_cond;
     n8_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue;
     n8_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output := n8_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1077_c2_8c24] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1077_c2_8c24] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1077_c2_8c24] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1077_c2_8c24] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output := result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1077_c2_8c24] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l1105_l1073_DUPLICATE_c0e4 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l1105_l1073_DUPLICATE_c0e4_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_04b4(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1077_c2_8c24_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l1105_l1073_DUPLICATE_c0e4_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l1105_l1073_DUPLICATE_c0e4_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
