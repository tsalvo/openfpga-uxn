-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity rot_0CLK_b288bfb7 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end rot_0CLK_b288bfb7;
architecture arch of rot_0CLK_b288bfb7 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal l8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_l8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2639_c6_35be]
signal BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2639_c2_8825]
signal result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2639_c2_8825]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2639_c2_8825]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2639_c2_8825]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2639_c2_8825]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2639_c2_8825]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2639_c2_8825]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2639_c2_8825]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2639_c2_8825]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2639_c2_8825]
signal l8_MUX_uxn_opcodes_h_l2639_c2_8825_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2639_c2_8825]
signal n8_MUX_uxn_opcodes_h_l2639_c2_8825_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2639_c2_8825]
signal t8_MUX_uxn_opcodes_h_l2639_c2_8825_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2652_c11_0cf2]
signal BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2652_c7_c8c2]
signal result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2652_c7_c8c2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2652_c7_c8c2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2652_c7_c8c2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2652_c7_c8c2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2652_c7_c8c2]
signal l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2652_c7_c8c2]
signal n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2652_c7_c8c2]
signal t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2655_c11_016a]
signal BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2655_c7_f145]
signal result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2655_c7_f145]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2655_c7_f145]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2655_c7_f145]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2655_c7_f145]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2655_c7_f145]
signal l8_MUX_uxn_opcodes_h_l2655_c7_f145_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2655_c7_f145_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2655_c7_f145]
signal n8_MUX_uxn_opcodes_h_l2655_c7_f145_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2655_c7_f145_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2655_c7_f145]
signal t8_MUX_uxn_opcodes_h_l2655_c7_f145_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2655_c7_f145_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2659_c11_ed3e]
signal BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2659_c7_33d3]
signal result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2659_c7_33d3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2659_c7_33d3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2659_c7_33d3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2659_c7_33d3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2659_c7_33d3]
signal l8_MUX_uxn_opcodes_h_l2659_c7_33d3_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2659_c7_33d3]
signal n8_MUX_uxn_opcodes_h_l2659_c7_33d3_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2661_c30_3fbd]
signal sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2666_c11_76db]
signal BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2666_c7_79d6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2666_c7_79d6]
signal result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2666_c7_79d6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2666_c7_79d6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2666_c7_79d6]
signal l8_MUX_uxn_opcodes_h_l2666_c7_79d6_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2672_c11_0503]
signal BIN_OP_EQ_uxn_opcodes_h_l2672_c11_0503_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2672_c11_0503_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2672_c11_0503_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2672_c7_462b]
signal result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2672_c7_462b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2672_c7_462b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_922a( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_vram_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_pc_updated := ref_toks_6;
      base.is_opc_done := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.is_stack_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be
BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_left,
BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_right,
BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_cond,
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_return_output);

-- l8_MUX_uxn_opcodes_h_l2639_c2_8825
l8_MUX_uxn_opcodes_h_l2639_c2_8825 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2639_c2_8825_cond,
l8_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue,
l8_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse,
l8_MUX_uxn_opcodes_h_l2639_c2_8825_return_output);

-- n8_MUX_uxn_opcodes_h_l2639_c2_8825
n8_MUX_uxn_opcodes_h_l2639_c2_8825 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2639_c2_8825_cond,
n8_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue,
n8_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse,
n8_MUX_uxn_opcodes_h_l2639_c2_8825_return_output);

-- t8_MUX_uxn_opcodes_h_l2639_c2_8825
t8_MUX_uxn_opcodes_h_l2639_c2_8825 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2639_c2_8825_cond,
t8_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue,
t8_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse,
t8_MUX_uxn_opcodes_h_l2639_c2_8825_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2
BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_left,
BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_right,
BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond,
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output);

-- l8_MUX_uxn_opcodes_h_l2652_c7_c8c2
l8_MUX_uxn_opcodes_h_l2652_c7_c8c2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond,
l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue,
l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse,
l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output);

-- n8_MUX_uxn_opcodes_h_l2652_c7_c8c2
n8_MUX_uxn_opcodes_h_l2652_c7_c8c2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond,
n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue,
n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse,
n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output);

-- t8_MUX_uxn_opcodes_h_l2652_c7_c8c2
t8_MUX_uxn_opcodes_h_l2652_c7_c8c2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond,
t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue,
t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse,
t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a
BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_left,
BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_right,
BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_cond,
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_return_output);

-- l8_MUX_uxn_opcodes_h_l2655_c7_f145
l8_MUX_uxn_opcodes_h_l2655_c7_f145 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2655_c7_f145_cond,
l8_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue,
l8_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse,
l8_MUX_uxn_opcodes_h_l2655_c7_f145_return_output);

-- n8_MUX_uxn_opcodes_h_l2655_c7_f145
n8_MUX_uxn_opcodes_h_l2655_c7_f145 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2655_c7_f145_cond,
n8_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue,
n8_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse,
n8_MUX_uxn_opcodes_h_l2655_c7_f145_return_output);

-- t8_MUX_uxn_opcodes_h_l2655_c7_f145
t8_MUX_uxn_opcodes_h_l2655_c7_f145 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2655_c7_f145_cond,
t8_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue,
t8_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse,
t8_MUX_uxn_opcodes_h_l2655_c7_f145_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e
BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_left,
BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_right,
BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_cond,
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output);

-- l8_MUX_uxn_opcodes_h_l2659_c7_33d3
l8_MUX_uxn_opcodes_h_l2659_c7_33d3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2659_c7_33d3_cond,
l8_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue,
l8_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse,
l8_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output);

-- n8_MUX_uxn_opcodes_h_l2659_c7_33d3
n8_MUX_uxn_opcodes_h_l2659_c7_33d3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2659_c7_33d3_cond,
n8_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue,
n8_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse,
n8_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd
sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_ins,
sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_x,
sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_y,
sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db
BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db_left,
BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db_right,
BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_cond,
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output);

-- l8_MUX_uxn_opcodes_h_l2666_c7_79d6
l8_MUX_uxn_opcodes_h_l2666_c7_79d6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2666_c7_79d6_cond,
l8_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue,
l8_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse,
l8_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2672_c11_0503
BIN_OP_EQ_uxn_opcodes_h_l2672_c11_0503 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2672_c11_0503_left,
BIN_OP_EQ_uxn_opcodes_h_l2672_c11_0503_right,
BIN_OP_EQ_uxn_opcodes_h_l2672_c11_0503_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_cond,
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 l8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_return_output,
 l8_MUX_uxn_opcodes_h_l2639_c2_8825_return_output,
 n8_MUX_uxn_opcodes_h_l2639_c2_8825_return_output,
 t8_MUX_uxn_opcodes_h_l2639_c2_8825_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output,
 l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output,
 n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output,
 t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_return_output,
 l8_MUX_uxn_opcodes_h_l2655_c7_f145_return_output,
 n8_MUX_uxn_opcodes_h_l2655_c7_f145_return_output,
 t8_MUX_uxn_opcodes_h_l2655_c7_f145_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output,
 l8_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output,
 n8_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output,
 sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output,
 l8_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2672_c11_0503_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2649_c3_45cb : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2644_c3_6999 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2639_c2_8825_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2639_c2_8825_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2639_c2_8825_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2639_c2_8825_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2653_c3_32da : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2655_c7_f145_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2655_c7_f145_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2655_c7_f145_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2656_c3_bac7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2655_c7_f145_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2655_c7_f145_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2655_c7_f145_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2663_c3_0354 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2659_c7_33d3_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2659_c7_33d3_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2668_c3_b360 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2669_c3_641b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2666_c7_79d6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_0503_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_0503_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_0503_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2673_c3_b69c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2672_c7_462b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2652_l2639_l2655_l2672_DUPLICATE_2add_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2652_l2666_l2655_DUPLICATE_1aa7_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2672_l2666_l2659_l2655_l2652_DUPLICATE_d6f9_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2659_l2652_l2655_DUPLICATE_16ac_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l2678_l2635_DUPLICATE_9788_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_l8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_l8 := l8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2656_c3_bac7 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2656_c3_bac7;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2673_c3_b69c := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2673_c3_b69c;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2649_c3_45cb := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2649_c3_45cb;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2663_c3_0354 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2663_c3_0354;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2653_c3_32da := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2653_c3_32da;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2668_c3_b360 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2668_c3_b360;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2644_c3_6999 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2644_c3_6999;
     VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_0503_right := to_unsigned(5, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2669_c3_641b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2669_c3_641b;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_ins := VAR_ins;
     VAR_l8_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse := l8;
     VAR_n8_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_0503_left := VAR_phase;
     VAR_l8_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse := t8;
     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2672_c7_462b] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2672_c7_462b_return_output := result.stack_address_sp_offset;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2639_c2_8825] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2639_c2_8825_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2659_l2652_l2655_DUPLICATE_16ac LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2659_l2652_l2655_DUPLICATE_16ac_return_output := result.is_stack_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2639_c2_8825] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2639_c2_8825_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l2666_c11_76db] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db_left;
     BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db_return_output := BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2639_c6_35be] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_left;
     BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_return_output := BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2652_c11_0cf2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_left;
     BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_return_output := BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2639_c2_8825] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2639_c2_8825_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2672_l2666_l2659_l2655_l2652_DUPLICATE_d6f9 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2672_l2666_l2659_l2655_l2652_DUPLICATE_d6f9_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2659_c11_ed3e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2652_l2639_l2655_l2672_DUPLICATE_2add LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2652_l2639_l2655_l2672_DUPLICATE_2add_return_output := result.u8_value;

     -- sp_relative_shift[uxn_opcodes_h_l2661_c30_3fbd] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_ins;
     sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_x;
     sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_return_output := sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2639_c2_8825] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2639_c2_8825_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2672_c11_0503] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2672_c11_0503_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_0503_left;
     BIN_OP_EQ_uxn_opcodes_h_l2672_c11_0503_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_0503_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_0503_return_output := BIN_OP_EQ_uxn_opcodes_h_l2672_c11_0503_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2652_l2666_l2655_DUPLICATE_1aa7 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2652_l2666_l2655_DUPLICATE_1aa7_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2655_c11_016a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_return_output;

     -- Submodule level 1
     VAR_l8_MUX_uxn_opcodes_h_l2639_c2_8825_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2639_c2_8825_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2639_c2_8825_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_35be_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_0cf2_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2655_c7_f145_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2655_c7_f145_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2655_c7_f145_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_016a_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2659_c7_33d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2659_c7_33d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_ed3e_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2666_c7_79d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_76db_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_0503_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_0503_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_0503_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2652_l2666_l2655_DUPLICATE_1aa7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2652_l2666_l2655_DUPLICATE_1aa7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2652_l2666_l2655_DUPLICATE_1aa7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2672_l2666_l2659_l2655_l2652_DUPLICATE_d6f9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2672_l2666_l2659_l2655_l2652_DUPLICATE_d6f9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2672_l2666_l2659_l2655_l2652_DUPLICATE_d6f9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2672_l2666_l2659_l2655_l2652_DUPLICATE_d6f9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2672_l2666_l2659_l2655_l2652_DUPLICATE_d6f9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2659_l2652_l2655_DUPLICATE_16ac_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2659_l2652_l2655_DUPLICATE_16ac_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2659_l2652_l2655_DUPLICATE_16ac_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2652_l2639_l2655_l2672_DUPLICATE_2add_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2652_l2639_l2655_l2672_DUPLICATE_2add_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2652_l2639_l2655_l2672_DUPLICATE_2add_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2652_l2639_l2655_l2672_DUPLICATE_2add_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2639_c2_8825_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2639_c2_8825_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2639_c2_8825_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2639_c2_8825_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2672_c7_462b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_3fbd_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2672_c7_462b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_return_output := result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2639_c2_8825] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2672_c7_462b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2639_c2_8825] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2672_c7_462b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2666_c7_79d6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output;

     -- t8_MUX[uxn_opcodes_h_l2655_c7_f145] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2655_c7_f145_cond <= VAR_t8_MUX_uxn_opcodes_h_l2655_c7_f145_cond;
     t8_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue;
     t8_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2655_c7_f145_return_output := t8_MUX_uxn_opcodes_h_l2655_c7_f145_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2639_c2_8825] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2659_c7_33d3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output;

     -- n8_MUX[uxn_opcodes_h_l2659_c7_33d3] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2659_c7_33d3_cond <= VAR_n8_MUX_uxn_opcodes_h_l2659_c7_33d3_cond;
     n8_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue;
     n8_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output := n8_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2639_c2_8825] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_return_output;

     -- l8_MUX[uxn_opcodes_h_l2666_c7_79d6] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2666_c7_79d6_cond <= VAR_l8_MUX_uxn_opcodes_h_l2666_c7_79d6_cond;
     l8_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue;
     l8_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output := l8_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output;

     -- Submodule level 2
     VAR_l8_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_462b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_462b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_462b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2655_c7_f145_return_output;
     -- l8_MUX[uxn_opcodes_h_l2659_c7_33d3] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2659_c7_33d3_cond <= VAR_l8_MUX_uxn_opcodes_h_l2659_c7_33d3_cond;
     l8_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue;
     l8_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output := l8_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output;

     -- t8_MUX[uxn_opcodes_h_l2652_c7_c8c2] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond <= VAR_t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond;
     t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue;
     t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output := t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2666_c7_79d6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output := result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2666_c7_79d6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output;

     -- n8_MUX[uxn_opcodes_h_l2655_c7_f145] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2655_c7_f145_cond <= VAR_n8_MUX_uxn_opcodes_h_l2655_c7_f145_cond;
     n8_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue;
     n8_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2655_c7_f145_return_output := n8_MUX_uxn_opcodes_h_l2655_c7_f145_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2666_c7_79d6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2655_c7_f145] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2659_c7_33d3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output;

     -- Submodule level 3
     VAR_l8_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2655_c7_f145_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_f145_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_79d6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output;
     -- l8_MUX[uxn_opcodes_h_l2655_c7_f145] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2655_c7_f145_cond <= VAR_l8_MUX_uxn_opcodes_h_l2655_c7_f145_cond;
     l8_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue;
     l8_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2655_c7_f145_return_output := l8_MUX_uxn_opcodes_h_l2655_c7_f145_return_output;

     -- t8_MUX[uxn_opcodes_h_l2639_c2_8825] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2639_c2_8825_cond <= VAR_t8_MUX_uxn_opcodes_h_l2639_c2_8825_cond;
     t8_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue;
     t8_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2639_c2_8825_return_output := t8_MUX_uxn_opcodes_h_l2639_c2_8825_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2659_c7_33d3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output := result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2659_c7_33d3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output;

     -- n8_MUX[uxn_opcodes_h_l2652_c7_c8c2] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond <= VAR_n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond;
     n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue;
     n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output := n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2659_c7_33d3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2652_c7_c8c2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2655_c7_f145] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_return_output;

     -- Submodule level 4
     VAR_l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2655_c7_f145_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_f145_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_33d3_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2639_c2_8825_return_output;
     -- l8_MUX[uxn_opcodes_h_l2652_c7_c8c2] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond <= VAR_l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond;
     l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue;
     l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output := l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2655_c7_f145] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_return_output := result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2639_c2_8825] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2652_c7_c8c2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2655_c7_f145] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2655_c7_f145] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_return_output;

     -- n8_MUX[uxn_opcodes_h_l2639_c2_8825] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2639_c2_8825_cond <= VAR_n8_MUX_uxn_opcodes_h_l2639_c2_8825_cond;
     n8_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue;
     n8_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2639_c2_8825_return_output := n8_MUX_uxn_opcodes_h_l2639_c2_8825_return_output;

     -- Submodule level 5
     VAR_l8_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output;
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2639_c2_8825_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_f145_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_f145_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_f145_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2652_c7_c8c2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2652_c7_c8c2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output := result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output;

     -- l8_MUX[uxn_opcodes_h_l2639_c2_8825] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2639_c2_8825_cond <= VAR_l8_MUX_uxn_opcodes_h_l2639_c2_8825_cond;
     l8_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue;
     l8_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2639_c2_8825_return_output := l8_MUX_uxn_opcodes_h_l2639_c2_8825_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2652_c7_c8c2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2639_c2_8825] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_return_output;

     -- Submodule level 6
     REG_VAR_l8 := VAR_l8_MUX_uxn_opcodes_h_l2639_c2_8825_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c8c2_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2639_c2_8825] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_return_output := result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2639_c2_8825] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2639_c2_8825] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l2678_l2635_DUPLICATE_9788 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l2678_l2635_DUPLICATE_9788_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_922a(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_8825_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_8825_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_8825_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_8825_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_8825_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_8825_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_8825_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_8825_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_8825_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l2678_l2635_DUPLICATE_9788_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l2678_l2635_DUPLICATE_9788_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_l8 <= REG_VAR_l8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     l8 <= REG_COMB_l8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
