-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 47
entity ldz_0CLK_b128164d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldz_0CLK_b128164d;
architecture arch of ldz_0CLK_b128164d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1437_c6_fb3c]
signal BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1437_c2_c008]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1437_c2_c008]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1437_c2_c008]
signal result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1437_c2_c008]
signal result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1437_c2_c008]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1437_c2_c008]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1437_c2_c008]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1437_c2_c008]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1437_c2_c008]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1437_c2_c008]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1437_c2_c008]
signal tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1437_c2_c008]
signal t8_MUX_uxn_opcodes_h_l1437_c2_c008_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1450_c11_68d5]
signal BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1450_c7_b34a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1450_c7_b34a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1450_c7_b34a]
signal result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1450_c7_b34a]
signal result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1450_c7_b34a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1450_c7_b34a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1450_c7_b34a]
signal tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1450_c7_b34a]
signal t8_MUX_uxn_opcodes_h_l1450_c7_b34a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1453_c11_deac]
signal BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1453_c7_943a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1453_c7_943a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1453_c7_943a]
signal result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1453_c7_943a]
signal result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1453_c7_943a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1453_c7_943a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1453_c7_943a]
signal tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1453_c7_943a]
signal t8_MUX_uxn_opcodes_h_l1453_c7_943a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1453_c7_943a_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1455_c30_4c0f]
signal sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1458_c11_50ef]
signal BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1458_c7_5df8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1458_c7_5df8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1458_c7_5df8]
signal result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1458_c7_5df8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1458_c7_5df8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1458_c7_5df8]
signal tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1461_c11_a25b]
signal BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1461_c7_0e34]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1461_c7_0e34]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1461_c7_0e34]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1461_c7_0e34]
signal result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1461_c7_0e34]
signal tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output : unsigned(7 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_500b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_pc_updated := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.u16_value := ref_toks_4;
      base.is_ram_write := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_stack_write := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_stack_index_flipped := ref_toks_9;
      base.is_opc_done := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c
BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_left,
BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_right,
BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008
result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008
result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008
result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_cond,
result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008
result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_cond,
result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008
result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1437_c2_c008
tmp8_MUX_uxn_opcodes_h_l1437_c2_c008 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_cond,
tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue,
tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse,
tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_return_output);

-- t8_MUX_uxn_opcodes_h_l1437_c2_c008
t8_MUX_uxn_opcodes_h_l1437_c2_c008 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1437_c2_c008_cond,
t8_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue,
t8_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse,
t8_MUX_uxn_opcodes_h_l1437_c2_c008_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5
BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_left,
BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_right,
BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a
result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a
result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_cond,
result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a
result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_cond,
result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a
tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_cond,
tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue,
tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse,
tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output);

-- t8_MUX_uxn_opcodes_h_l1450_c7_b34a
t8_MUX_uxn_opcodes_h_l1450_c7_b34a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1450_c7_b34a_cond,
t8_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue,
t8_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse,
t8_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac
BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_left,
BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_right,
BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a
result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a
result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a
result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_cond,
result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a
result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_cond,
result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a
result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1453_c7_943a
tmp8_MUX_uxn_opcodes_h_l1453_c7_943a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_cond,
tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue,
tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse,
tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_return_output);

-- t8_MUX_uxn_opcodes_h_l1453_c7_943a
t8_MUX_uxn_opcodes_h_l1453_c7_943a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1453_c7_943a_cond,
t8_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue,
t8_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse,
t8_MUX_uxn_opcodes_h_l1453_c7_943a_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f
sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_ins,
sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_x,
sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_y,
sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef
BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef_left,
BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef_right,
BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8
result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8
result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8
result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_cond,
result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8
result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8
tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_cond,
tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue,
tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse,
tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b
BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b_left,
BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b_right,
BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34
result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34
result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34
result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_cond,
result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34
tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_cond,
tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue,
tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse,
tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_return_output,
 tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_return_output,
 t8_MUX_uxn_opcodes_h_l1437_c2_c008_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output,
 tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output,
 t8_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_return_output,
 tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_return_output,
 t8_MUX_uxn_opcodes_h_l1453_c7_943a_return_output,
 sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output,
 tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output,
 tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1442_c3_8fed : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1447_c3_bb41 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1437_c2_c008_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1437_c2_c008_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1451_c3_a928 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1453_c7_943a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1450_c7_b34a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1453_c7_943a_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1456_c22_ba5a_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1459_c3_47c8 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1464_c3_23dc : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1461_l1458_l1453_l1450_l1437_DUPLICATE_cfb1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1437_l1450_l1453_DUPLICATE_184f_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1458_l1450_DUPLICATE_9a19_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_0558_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_8456_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1458_l1461_l1453_DUPLICATE_53bb_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_500b_uxn_opcodes_h_l1469_l1433_DUPLICATE_88f5_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1447_c3_bb41 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1447_c3_bb41;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1464_c3_23dc := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1464_c3_23dc;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1451_c3_a928 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1451_c3_a928;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_right := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1459_c3_47c8 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1459_c3_47c8;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1442_c3_8fed := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1442_c3_8fed;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b_right := to_unsigned(4, 3);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse := tmp8;
     -- sp_relative_shift[uxn_opcodes_h_l1455_c30_4c0f] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_ins;
     sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_x;
     sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_return_output := sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1437_c2_c008] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1437_c2_c008_return_output := result.is_pc_updated;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1437_c2_c008] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1437_c2_c008_return_output := result.is_ram_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1437_c2_c008] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1437_c2_c008_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1458_l1450_DUPLICATE_9a19 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1458_l1450_DUPLICATE_9a19_return_output := result.sp_relative_shift;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1456_c22_ba5a] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1456_c22_ba5a_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1437_l1450_l1453_DUPLICATE_184f LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1437_l1450_l1453_DUPLICATE_184f_return_output := result.u16_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1453_c11_deac] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_left;
     BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_return_output := BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1461_l1458_l1453_l1450_l1437_DUPLICATE_cfb1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1461_l1458_l1453_l1450_l1437_DUPLICATE_cfb1_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1461_c11_a25b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_0558 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_0558_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1437_c6_fb3c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1450_c11_68d5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_left;
     BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_return_output := BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1458_c11_50ef] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef_left;
     BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef_return_output := BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1437_c2_c008] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1437_c2_c008_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1458_l1461_l1453_DUPLICATE_53bb LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1458_l1461_l1453_DUPLICATE_53bb_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_8456 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_8456_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1437_c2_c008_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_fb3c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1450_c7_b34a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_68d5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1453_c7_943a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_deac_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_50ef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_a25b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1456_c22_ba5a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1458_l1450_DUPLICATE_9a19_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1458_l1450_DUPLICATE_9a19_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1437_l1450_l1453_DUPLICATE_184f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1437_l1450_l1453_DUPLICATE_184f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1437_l1450_l1453_DUPLICATE_184f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_8456_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_8456_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_8456_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_8456_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_0558_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_0558_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_0558_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_0558_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1458_l1461_l1453_DUPLICATE_53bb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1458_l1461_l1453_DUPLICATE_53bb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1458_l1461_l1453_DUPLICATE_53bb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1461_l1458_l1453_l1450_l1437_DUPLICATE_cfb1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1461_l1458_l1453_l1450_l1437_DUPLICATE_cfb1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1461_l1458_l1453_l1450_l1437_DUPLICATE_cfb1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1461_l1458_l1453_l1450_l1437_DUPLICATE_cfb1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1461_l1458_l1453_l1450_l1437_DUPLICATE_cfb1_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1437_c2_c008_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1437_c2_c008_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1437_c2_c008_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1437_c2_c008_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_4c0f_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1461_c7_0e34] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output := result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1461_c7_0e34] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1437_c2_c008] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1461_c7_0e34] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1458_c7_5df8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1437_c2_c008] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1453_c7_943a] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_return_output := result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1461_c7_0e34] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1437_c2_c008] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_return_output;

     -- t8_MUX[uxn_opcodes_h_l1453_c7_943a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1453_c7_943a_cond <= VAR_t8_MUX_uxn_opcodes_h_l1453_c7_943a_cond;
     t8_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue;
     t8_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1453_c7_943a_return_output := t8_MUX_uxn_opcodes_h_l1453_c7_943a_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1461_c7_0e34] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_cond;
     tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output := tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1437_c2_c008] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_943a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1453_c7_943a_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_0e34_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1458_c7_5df8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output := result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1458_c7_5df8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1458_c7_5df8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output;

     -- t8_MUX[uxn_opcodes_h_l1450_c7_b34a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1450_c7_b34a_cond <= VAR_t8_MUX_uxn_opcodes_h_l1450_c7_b34a_cond;
     t8_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue;
     t8_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output := t8_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1453_c7_943a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1450_c7_b34a] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output := result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1458_c7_5df8] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_cond;
     tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output := tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1458_c7_5df8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_943a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_5df8_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1453_c7_943a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1453_c7_943a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_return_output := result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1450_c7_b34a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1453_c7_943a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1437_c2_c008] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_return_output := result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1453_c7_943a] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_cond;
     tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_return_output := tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1453_c7_943a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_return_output;

     -- t8_MUX[uxn_opcodes_h_l1437_c2_c008] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1437_c2_c008_cond <= VAR_t8_MUX_uxn_opcodes_h_l1437_c2_c008_cond;
     t8_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue;
     t8_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1437_c2_c008_return_output := t8_MUX_uxn_opcodes_h_l1437_c2_c008_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_943a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_943a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_943a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_943a_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1437_c2_c008_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_943a_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1450_c7_b34a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output := result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1437_c2_c008] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1450_c7_b34a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1450_c7_b34a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1450_c7_b34a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1450_c7_b34a] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_cond;
     tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output := tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_b34a_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1437_c2_c008] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1437_c2_c008] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1437_c2_c008] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1437_c2_c008] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_return_output := result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1437_c2_c008] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_cond;
     tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_return_output := tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_return_output;

     -- Submodule level 6
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_c008_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_500b_uxn_opcodes_h_l1469_l1433_DUPLICATE_88f5 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_500b_uxn_opcodes_h_l1469_l1433_DUPLICATE_88f5_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_500b(
     result,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_c008_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_c008_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_c008_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_c008_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_c008_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_c008_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_c008_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_c008_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_c008_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_c008_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_500b_uxn_opcodes_h_l1469_l1433_DUPLICATE_88f5_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_500b_uxn_opcodes_h_l1469_l1433_DUPLICATE_88f5_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
