-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity lth_0CLK_85d5529e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end lth_0CLK_85d5529e;
architecture arch of lth_0CLK_85d5529e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1800_c6_4525]
signal BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1800_c1_b4d4]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1800_c2_5caa]
signal n8_MUX_uxn_opcodes_h_l1800_c2_5caa_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1800_c2_5caa]
signal t8_MUX_uxn_opcodes_h_l1800_c2_5caa_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1800_c2_5caa]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1800_c2_5caa]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1800_c2_5caa]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1800_c2_5caa]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1800_c2_5caa]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1800_c2_5caa]
signal result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1801_c3_5c7f[uxn_opcodes_h_l1801_c3_5c7f]
signal printf_uxn_opcodes_h_l1801_c3_5c7f_uxn_opcodes_h_l1801_c3_5c7f_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1805_c11_a1d8]
signal BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1805_c7_2076]
signal n8_MUX_uxn_opcodes_h_l1805_c7_2076_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1805_c7_2076_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1805_c7_2076]
signal t8_MUX_uxn_opcodes_h_l1805_c7_2076_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1805_c7_2076_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1805_c7_2076]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1805_c7_2076]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1805_c7_2076]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1805_c7_2076]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1805_c7_2076]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1805_c7_2076]
signal result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1808_c11_0402]
signal BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1808_c7_b315]
signal n8_MUX_uxn_opcodes_h_l1808_c7_b315_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1808_c7_b315_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1808_c7_b315]
signal t8_MUX_uxn_opcodes_h_l1808_c7_b315_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1808_c7_b315_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1808_c7_b315]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1808_c7_b315]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1808_c7_b315]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1808_c7_b315]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1808_c7_b315]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1808_c7_b315]
signal result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1811_c11_095a]
signal BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1811_c7_7003]
signal n8_MUX_uxn_opcodes_h_l1811_c7_7003_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1811_c7_7003_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1811_c7_7003]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1811_c7_7003]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1811_c7_7003]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1811_c7_7003]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1811_c7_7003]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1811_c7_7003]
signal result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1814_c30_7c7f]
signal sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_return_output : signed(3 downto 0);

-- BIN_OP_LT[uxn_opcodes_h_l1817_c21_472f]
signal BIN_OP_LT_uxn_opcodes_h_l1817_c21_472f_left : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l1817_c21_472f_right : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l1817_c21_472f_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1817_c21_1618]
signal MUX_uxn_opcodes_h_l1817_c21_1618_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1817_c21_1618_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1817_c21_1618_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1817_c21_1618_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1819_c11_ef0c]
signal BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ef0c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ef0c_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ef0c_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1819_c7_acb4]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1819_c7_acb4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1819_c7_acb4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_5b93( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525
BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_left,
BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_right,
BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_return_output);

-- n8_MUX_uxn_opcodes_h_l1800_c2_5caa
n8_MUX_uxn_opcodes_h_l1800_c2_5caa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1800_c2_5caa_cond,
n8_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue,
n8_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse,
n8_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output);

-- t8_MUX_uxn_opcodes_h_l1800_c2_5caa
t8_MUX_uxn_opcodes_h_l1800_c2_5caa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1800_c2_5caa_cond,
t8_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue,
t8_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse,
t8_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa
result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa
result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa
result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa
result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa
result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_cond,
result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output);

-- printf_uxn_opcodes_h_l1801_c3_5c7f_uxn_opcodes_h_l1801_c3_5c7f
printf_uxn_opcodes_h_l1801_c3_5c7f_uxn_opcodes_h_l1801_c3_5c7f : entity work.printf_uxn_opcodes_h_l1801_c3_5c7f_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1801_c3_5c7f_uxn_opcodes_h_l1801_c3_5c7f_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8
BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_left,
BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_right,
BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_return_output);

-- n8_MUX_uxn_opcodes_h_l1805_c7_2076
n8_MUX_uxn_opcodes_h_l1805_c7_2076 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1805_c7_2076_cond,
n8_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue,
n8_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse,
n8_MUX_uxn_opcodes_h_l1805_c7_2076_return_output);

-- t8_MUX_uxn_opcodes_h_l1805_c7_2076
t8_MUX_uxn_opcodes_h_l1805_c7_2076 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1805_c7_2076_cond,
t8_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue,
t8_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse,
t8_MUX_uxn_opcodes_h_l1805_c7_2076_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076
result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076
result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076
result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076
result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076
result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_cond,
result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402
BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_left,
BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_right,
BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_return_output);

-- n8_MUX_uxn_opcodes_h_l1808_c7_b315
n8_MUX_uxn_opcodes_h_l1808_c7_b315 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1808_c7_b315_cond,
n8_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue,
n8_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse,
n8_MUX_uxn_opcodes_h_l1808_c7_b315_return_output);

-- t8_MUX_uxn_opcodes_h_l1808_c7_b315
t8_MUX_uxn_opcodes_h_l1808_c7_b315 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1808_c7_b315_cond,
t8_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue,
t8_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse,
t8_MUX_uxn_opcodes_h_l1808_c7_b315_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315
result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315
result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315
result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315
result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315
result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_cond,
result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a
BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_left,
BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_right,
BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_return_output);

-- n8_MUX_uxn_opcodes_h_l1811_c7_7003
n8_MUX_uxn_opcodes_h_l1811_c7_7003 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1811_c7_7003_cond,
n8_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue,
n8_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse,
n8_MUX_uxn_opcodes_h_l1811_c7_7003_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003
result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003
result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003
result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003
result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003
result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_cond,
result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f
sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_ins,
sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_x,
sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_y,
sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_return_output);

-- BIN_OP_LT_uxn_opcodes_h_l1817_c21_472f
BIN_OP_LT_uxn_opcodes_h_l1817_c21_472f : entity work.BIN_OP_LT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_LT_uxn_opcodes_h_l1817_c21_472f_left,
BIN_OP_LT_uxn_opcodes_h_l1817_c21_472f_right,
BIN_OP_LT_uxn_opcodes_h_l1817_c21_472f_return_output);

-- MUX_uxn_opcodes_h_l1817_c21_1618
MUX_uxn_opcodes_h_l1817_c21_1618 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1817_c21_1618_cond,
MUX_uxn_opcodes_h_l1817_c21_1618_iftrue,
MUX_uxn_opcodes_h_l1817_c21_1618_iffalse,
MUX_uxn_opcodes_h_l1817_c21_1618_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ef0c
BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ef0c : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ef0c_left,
BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ef0c_right,
BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ef0c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4
result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4
result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4
result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_return_output,
 n8_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output,
 t8_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_return_output,
 n8_MUX_uxn_opcodes_h_l1805_c7_2076_return_output,
 t8_MUX_uxn_opcodes_h_l1805_c7_2076_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_return_output,
 n8_MUX_uxn_opcodes_h_l1808_c7_b315_return_output,
 t8_MUX_uxn_opcodes_h_l1808_c7_b315_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_return_output,
 n8_MUX_uxn_opcodes_h_l1811_c7_7003_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_return_output,
 sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_return_output,
 BIN_OP_LT_uxn_opcodes_h_l1817_c21_472f_return_output,
 MUX_uxn_opcodes_h_l1817_c21_1618_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ef0c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1805_c7_2076_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1800_c2_5caa_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1805_c7_2076_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1800_c2_5caa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1802_c3_de53 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1801_c3_5c7f_uxn_opcodes_h_l1801_c3_5c7f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1808_c7_b315_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1805_c7_2076_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1808_c7_b315_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1805_c7_2076_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1806_c3_55e5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1811_c7_7003_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1808_c7_b315_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1808_c7_b315_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1811_c7_7003_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1816_c3_3475 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1817_c21_1618_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1817_c21_1618_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1817_c21_1618_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_472f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_472f_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_472f_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1817_c21_1618_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ef0c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ef0c_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ef0c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1800_l1805_l1819_l1808_DUPLICATE_64ba_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1800_l1805_l1819_l1808_DUPLICATE_3819_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1800_l1811_l1805_l1808_DUPLICATE_f615_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1800_l1811_l1805_l1808_DUPLICATE_70dc_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1811_l1805_l1819_l1808_DUPLICATE_a458_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1811_l1808_DUPLICATE_1fda_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1825_l1796_DUPLICATE_7ba0_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1806_c3_55e5 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1806_c3_55e5;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ef0c_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1802_c3_de53 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1802_c3_de53;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_iffalse := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1817_c21_1618_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1817_c21_1618_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1816_c3_3475 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1816_c3_3475;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ef0c_left := VAR_phase;
     VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_472f_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_472f_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse := t8;
     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1800_l1811_l1805_l1808_DUPLICATE_70dc LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1800_l1811_l1805_l1808_DUPLICATE_70dc_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1800_c6_4525] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_left;
     BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_return_output := BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1808_c11_0402] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_left;
     BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_return_output := BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_return_output;

     -- BIN_OP_LT[uxn_opcodes_h_l1817_c21_472f] LATENCY=0
     -- Inputs
     BIN_OP_LT_uxn_opcodes_h_l1817_c21_472f_left <= VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_472f_left;
     BIN_OP_LT_uxn_opcodes_h_l1817_c21_472f_right <= VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_472f_right;
     -- Outputs
     VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_472f_return_output := BIN_OP_LT_uxn_opcodes_h_l1817_c21_472f_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1800_l1805_l1819_l1808_DUPLICATE_3819 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1800_l1805_l1819_l1808_DUPLICATE_3819_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1819_c11_ef0c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ef0c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ef0c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ef0c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ef0c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ef0c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ef0c_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1814_c30_7c7f] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_ins;
     sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_x;
     sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_return_output := sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1800_l1805_l1819_l1808_DUPLICATE_64ba LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1800_l1805_l1819_l1808_DUPLICATE_64ba_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1805_c11_a1d8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_left;
     BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_return_output := BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1811_c11_095a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1811_l1805_l1819_l1808_DUPLICATE_a458 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1811_l1805_l1819_l1808_DUPLICATE_a458_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1811_l1808_DUPLICATE_1fda LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1811_l1808_DUPLICATE_1fda_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1800_l1811_l1805_l1808_DUPLICATE_f615 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1800_l1811_l1805_l1808_DUPLICATE_f615_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1800_c2_5caa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1800_c2_5caa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_4525_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1805_c7_2076_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1805_c7_2076_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_a1d8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1808_c7_b315_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1808_c7_b315_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_0402_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1811_c7_7003_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_095a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ef0c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ef0c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ef0c_return_output;
     VAR_MUX_uxn_opcodes_h_l1817_c21_1618_cond := VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_472f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1800_l1811_l1805_l1808_DUPLICATE_f615_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1800_l1811_l1805_l1808_DUPLICATE_f615_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1800_l1811_l1805_l1808_DUPLICATE_f615_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1800_l1811_l1805_l1808_DUPLICATE_f615_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1811_l1805_l1819_l1808_DUPLICATE_a458_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1811_l1805_l1819_l1808_DUPLICATE_a458_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1811_l1805_l1819_l1808_DUPLICATE_a458_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1811_l1805_l1819_l1808_DUPLICATE_a458_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1800_l1805_l1819_l1808_DUPLICATE_3819_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1800_l1805_l1819_l1808_DUPLICATE_3819_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1800_l1805_l1819_l1808_DUPLICATE_3819_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1800_l1805_l1819_l1808_DUPLICATE_3819_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1800_l1805_l1819_l1808_DUPLICATE_64ba_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1800_l1805_l1819_l1808_DUPLICATE_64ba_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1800_l1805_l1819_l1808_DUPLICATE_64ba_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1800_l1805_l1819_l1808_DUPLICATE_64ba_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1811_l1808_DUPLICATE_1fda_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1811_l1808_DUPLICATE_1fda_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1800_l1811_l1805_l1808_DUPLICATE_70dc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1800_l1811_l1805_l1808_DUPLICATE_70dc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1800_l1811_l1805_l1808_DUPLICATE_70dc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1800_l1811_l1805_l1808_DUPLICATE_70dc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_7c7f_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1811_c7_7003] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1811_c7_7003] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1819_c7_acb4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_return_output;

     -- n8_MUX[uxn_opcodes_h_l1811_c7_7003] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1811_c7_7003_cond <= VAR_n8_MUX_uxn_opcodes_h_l1811_c7_7003_cond;
     n8_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue;
     n8_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1811_c7_7003_return_output := n8_MUX_uxn_opcodes_h_l1811_c7_7003_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1819_c7_acb4] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1819_c7_acb4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_return_output;

     -- t8_MUX[uxn_opcodes_h_l1808_c7_b315] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1808_c7_b315_cond <= VAR_t8_MUX_uxn_opcodes_h_l1808_c7_b315_cond;
     t8_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue;
     t8_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1808_c7_b315_return_output := t8_MUX_uxn_opcodes_h_l1808_c7_b315_return_output;

     -- MUX[uxn_opcodes_h_l1817_c21_1618] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1817_c21_1618_cond <= VAR_MUX_uxn_opcodes_h_l1817_c21_1618_cond;
     MUX_uxn_opcodes_h_l1817_c21_1618_iftrue <= VAR_MUX_uxn_opcodes_h_l1817_c21_1618_iftrue;
     MUX_uxn_opcodes_h_l1817_c21_1618_iffalse <= VAR_MUX_uxn_opcodes_h_l1817_c21_1618_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1817_c21_1618_return_output := MUX_uxn_opcodes_h_l1817_c21_1618_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1800_c1_b4d4] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue := VAR_MUX_uxn_opcodes_h_l1817_c21_1618_return_output;
     VAR_printf_uxn_opcodes_h_l1801_c3_5c7f_uxn_opcodes_h_l1801_c3_5c7f_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_b4d4_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1811_c7_7003_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_acb4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_acb4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_acb4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7003_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7003_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1808_c7_b315_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1811_c7_7003] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1811_c7_7003] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_return_output := result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_return_output;

     -- t8_MUX[uxn_opcodes_h_l1805_c7_2076] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1805_c7_2076_cond <= VAR_t8_MUX_uxn_opcodes_h_l1805_c7_2076_cond;
     t8_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue;
     t8_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1805_c7_2076_return_output := t8_MUX_uxn_opcodes_h_l1805_c7_2076_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1808_c7_b315] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_return_output;

     -- printf_uxn_opcodes_h_l1801_c3_5c7f[uxn_opcodes_h_l1801_c3_5c7f] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1801_c3_5c7f_uxn_opcodes_h_l1801_c3_5c7f_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1801_c3_5c7f_uxn_opcodes_h_l1801_c3_5c7f_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1811_c7_7003] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_return_output;

     -- n8_MUX[uxn_opcodes_h_l1808_c7_b315] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1808_c7_b315_cond <= VAR_n8_MUX_uxn_opcodes_h_l1808_c7_b315_cond;
     n8_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue;
     n8_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1808_c7_b315_return_output := n8_MUX_uxn_opcodes_h_l1808_c7_b315_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1808_c7_b315] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1811_c7_7003] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1808_c7_b315_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7003_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7003_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7003_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_b315_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_b315_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7003_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1805_c7_2076_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1808_c7_b315] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_return_output;

     -- n8_MUX[uxn_opcodes_h_l1805_c7_2076] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1805_c7_2076_cond <= VAR_n8_MUX_uxn_opcodes_h_l1805_c7_2076_cond;
     n8_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue;
     n8_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1805_c7_2076_return_output := n8_MUX_uxn_opcodes_h_l1805_c7_2076_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1808_c7_b315] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1805_c7_2076] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_return_output;

     -- t8_MUX[uxn_opcodes_h_l1800_c2_5caa] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1800_c2_5caa_cond <= VAR_t8_MUX_uxn_opcodes_h_l1800_c2_5caa_cond;
     t8_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue;
     t8_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output := t8_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1808_c7_b315] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_return_output := result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1808_c7_b315] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1805_c7_2076] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1805_c7_2076_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_b315_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_b315_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_b315_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_2076_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_2076_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_b315_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1805_c7_2076] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1805_c7_2076] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_return_output := result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1805_c7_2076] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_return_output;

     -- n8_MUX[uxn_opcodes_h_l1800_c2_5caa] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1800_c2_5caa_cond <= VAR_n8_MUX_uxn_opcodes_h_l1800_c2_5caa_cond;
     n8_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue;
     n8_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output := n8_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1800_c2_5caa] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1805_c7_2076] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1800_c2_5caa] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_2076_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_2076_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_2076_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_2076_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1800_c2_5caa] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output := result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1800_c2_5caa] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1800_c2_5caa] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1800_c2_5caa] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1825_l1796_DUPLICATE_7ba0 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1825_l1796_DUPLICATE_7ba0_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5b93(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_5caa_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1825_l1796_DUPLICATE_7ba0_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1825_l1796_DUPLICATE_7ba0_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
