-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity div_0CLK_4e24eea7 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end div_0CLK_4e24eea7;
architecture arch of div_0CLK_4e24eea7 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2056_c6_3787]
signal BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2056_c2_5cb8]
signal n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2056_c2_5cb8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2056_c2_5cb8]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2056_c2_5cb8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2056_c2_5cb8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2056_c2_5cb8]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2056_c2_5cb8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2056_c2_5cb8]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2056_c2_5cb8]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2056_c2_5cb8]
signal result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2056_c2_5cb8]
signal t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2069_c11_6e4f]
signal BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2069_c7_fea5]
signal n8_MUX_uxn_opcodes_h_l2069_c7_fea5_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2069_c7_fea5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2069_c7_fea5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2069_c7_fea5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2069_c7_fea5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2069_c7_fea5]
signal result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2069_c7_fea5]
signal t8_MUX_uxn_opcodes_h_l2069_c7_fea5_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2072_c11_4c96]
signal BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2072_c7_d6ad]
signal n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2072_c7_d6ad]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2072_c7_d6ad]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2072_c7_d6ad]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2072_c7_d6ad]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2072_c7_d6ad]
signal result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2072_c7_d6ad]
signal t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2075_c11_91f0]
signal BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2075_c7_71b6]
signal n8_MUX_uxn_opcodes_h_l2075_c7_71b6_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2075_c7_71b6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2075_c7_71b6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2075_c7_71b6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2075_c7_71b6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2075_c7_71b6]
signal result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2077_c30_f128]
signal sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2080_c21_6cca]
signal BIN_OP_EQ_uxn_opcodes_h_l2080_c21_6cca_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2080_c21_6cca_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2080_c21_6cca_return_output : unsigned(0 downto 0);

-- BIN_OP_DIV[uxn_opcodes_h_l2080_c35_93a1]
signal BIN_OP_DIV_uxn_opcodes_h_l2080_c35_93a1_left : unsigned(7 downto 0);
signal BIN_OP_DIV_uxn_opcodes_h_l2080_c35_93a1_right : unsigned(7 downto 0);
signal BIN_OP_DIV_uxn_opcodes_h_l2080_c35_93a1_return_output : unsigned(7 downto 0);

-- MUX[uxn_opcodes_h_l2080_c21_ce84]
signal MUX_uxn_opcodes_h_l2080_c21_ce84_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l2080_c21_ce84_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l2080_c21_ce84_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l2080_c21_ce84_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_04b4( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.is_stack_index_flipped := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.u8_value := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787
BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_left,
BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_right,
BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_return_output);

-- n8_MUX_uxn_opcodes_h_l2056_c2_5cb8
n8_MUX_uxn_opcodes_h_l2056_c2_5cb8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond,
n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue,
n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse,
n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8
result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8
result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8
result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8
result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8
result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8
result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8
result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond,
result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output);

-- t8_MUX_uxn_opcodes_h_l2056_c2_5cb8
t8_MUX_uxn_opcodes_h_l2056_c2_5cb8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond,
t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue,
t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse,
t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f
BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_left,
BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_right,
BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_return_output);

-- n8_MUX_uxn_opcodes_h_l2069_c7_fea5
n8_MUX_uxn_opcodes_h_l2069_c7_fea5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2069_c7_fea5_cond,
n8_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue,
n8_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse,
n8_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5
result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5
result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5
result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5
result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_cond,
result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output);

-- t8_MUX_uxn_opcodes_h_l2069_c7_fea5
t8_MUX_uxn_opcodes_h_l2069_c7_fea5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2069_c7_fea5_cond,
t8_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue,
t8_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse,
t8_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96
BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_left,
BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_right,
BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_return_output);

-- n8_MUX_uxn_opcodes_h_l2072_c7_d6ad
n8_MUX_uxn_opcodes_h_l2072_c7_d6ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond,
n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue,
n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse,
n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad
result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad
result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad
result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad
result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond,
result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output);

-- t8_MUX_uxn_opcodes_h_l2072_c7_d6ad
t8_MUX_uxn_opcodes_h_l2072_c7_d6ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond,
t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue,
t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse,
t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0
BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0_left,
BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0_right,
BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0_return_output);

-- n8_MUX_uxn_opcodes_h_l2075_c7_71b6
n8_MUX_uxn_opcodes_h_l2075_c7_71b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2075_c7_71b6_cond,
n8_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue,
n8_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse,
n8_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6
result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6
result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6
result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6
result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_cond,
result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2077_c30_f128
sp_relative_shift_uxn_opcodes_h_l2077_c30_f128 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_ins,
sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_x,
sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_y,
sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2080_c21_6cca
BIN_OP_EQ_uxn_opcodes_h_l2080_c21_6cca : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2080_c21_6cca_left,
BIN_OP_EQ_uxn_opcodes_h_l2080_c21_6cca_right,
BIN_OP_EQ_uxn_opcodes_h_l2080_c21_6cca_return_output);

-- BIN_OP_DIV_uxn_opcodes_h_l2080_c35_93a1
BIN_OP_DIV_uxn_opcodes_h_l2080_c35_93a1 : entity work.BIN_OP_DIV_uint8_t_uint8_t_0CLK_371b3c10 port map (
BIN_OP_DIV_uxn_opcodes_h_l2080_c35_93a1_left,
BIN_OP_DIV_uxn_opcodes_h_l2080_c35_93a1_right,
BIN_OP_DIV_uxn_opcodes_h_l2080_c35_93a1_return_output);

-- MUX_uxn_opcodes_h_l2080_c21_ce84
MUX_uxn_opcodes_h_l2080_c21_ce84 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l2080_c21_ce84_cond,
MUX_uxn_opcodes_h_l2080_c21_ce84_iftrue,
MUX_uxn_opcodes_h_l2080_c21_ce84_iffalse,
MUX_uxn_opcodes_h_l2080_c21_ce84_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_return_output,
 n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output,
 t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_return_output,
 n8_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output,
 t8_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_return_output,
 n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output,
 t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0_return_output,
 n8_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output,
 sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2080_c21_6cca_return_output,
 BIN_OP_DIV_uxn_opcodes_h_l2080_c35_93a1_return_output,
 MUX_uxn_opcodes_h_l2080_c21_ce84_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2056_c2_5cb8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2066_c3_1718 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2056_c2_5cb8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2061_c3_5478 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2056_c2_5cb8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2056_c2_5cb8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2069_c7_fea5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2070_c3_ddae : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2069_c7_fea5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2075_c7_71b6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2079_c3_ccf9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2080_c21_ce84_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_6cca_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_6cca_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_6cca_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2080_c21_ce84_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2080_c21_ce84_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_93a1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_93a1_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_93a1_return_output : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2080_c21_ce84_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2069_l2072_l2056_l2075_DUPLICATE_e957_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2069_l2072_l2075_DUPLICATE_aece_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2069_l2072_l2075_DUPLICATE_7ec2_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2069_l2072_l2075_DUPLICATE_27fa_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2072_l2075_DUPLICATE_6ce0_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2052_l2084_DUPLICATE_574d_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2066_c3_1718 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2066_c3_1718;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l2080_c21_ce84_iftrue := resize(to_unsigned(0, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2079_c3_ccf9 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2079_c3_ccf9;
     VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_6cca_right := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2061_c3_5478 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2061_c3_5478;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2070_c3_ddae := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2070_c3_ddae;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_right := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0_left := VAR_phase;
     VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_93a1_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_93a1_right := t8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_6cca_left := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2069_l2072_l2075_DUPLICATE_7ec2 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2069_l2072_l2075_DUPLICATE_7ec2_return_output := result.is_opc_done;

     -- sp_relative_shift[uxn_opcodes_h_l2077_c30_f128] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_ins;
     sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_x;
     sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_return_output := sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2056_c2_5cb8] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2056_c2_5cb8_return_output := result.is_ram_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2069_l2072_l2075_DUPLICATE_aece LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2069_l2072_l2075_DUPLICATE_aece_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2069_c11_6e4f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_return_output;

     -- BIN_OP_DIV[uxn_opcodes_h_l2080_c35_93a1] LATENCY=0
     -- Inputs
     BIN_OP_DIV_uxn_opcodes_h_l2080_c35_93a1_left <= VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_93a1_left;
     BIN_OP_DIV_uxn_opcodes_h_l2080_c35_93a1_right <= VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_93a1_right;
     -- Outputs
     VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_93a1_return_output := BIN_OP_DIV_uxn_opcodes_h_l2080_c35_93a1_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2069_l2072_l2056_l2075_DUPLICATE_e957 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2069_l2072_l2056_l2075_DUPLICATE_e957_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2080_c21_6cca] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2080_c21_6cca_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_6cca_left;
     BIN_OP_EQ_uxn_opcodes_h_l2080_c21_6cca_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_6cca_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_6cca_return_output := BIN_OP_EQ_uxn_opcodes_h_l2080_c21_6cca_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2056_c2_5cb8] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2056_c2_5cb8_return_output := result.is_vram_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2056_c2_5cb8] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2056_c2_5cb8_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l2075_c11_91f0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0_left;
     BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0_return_output := BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2056_c6_3787] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_left;
     BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_return_output := BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2072_c11_4c96] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_left;
     BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_return_output := BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2072_l2075_DUPLICATE_6ce0 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2072_l2075_DUPLICATE_6ce0_return_output := result.stack_address_sp_offset;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2056_c2_5cb8] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2056_c2_5cb8_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2069_l2072_l2075_DUPLICATE_27fa LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2069_l2072_l2075_DUPLICATE_27fa_return_output := result.is_stack_write;

     -- Submodule level 1
     VAR_MUX_uxn_opcodes_h_l2080_c21_ce84_iffalse := VAR_BIN_OP_DIV_uxn_opcodes_h_l2080_c35_93a1_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2056_c6_3787_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2069_c7_fea5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2069_c7_fea5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_6e4f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2072_c11_4c96_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2075_c7_71b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2075_c11_91f0_return_output;
     VAR_MUX_uxn_opcodes_h_l2080_c21_ce84_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2080_c21_6cca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2069_l2072_l2075_DUPLICATE_aece_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2069_l2072_l2075_DUPLICATE_aece_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2069_l2072_l2075_DUPLICATE_aece_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2069_l2072_l2075_DUPLICATE_7ec2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2069_l2072_l2075_DUPLICATE_7ec2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2069_l2072_l2075_DUPLICATE_7ec2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2069_l2072_l2075_DUPLICATE_27fa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2069_l2072_l2075_DUPLICATE_27fa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2069_l2072_l2075_DUPLICATE_27fa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2072_l2075_DUPLICATE_6ce0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2072_l2075_DUPLICATE_6ce0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2069_l2072_l2056_l2075_DUPLICATE_e957_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2069_l2072_l2056_l2075_DUPLICATE_e957_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2069_l2072_l2056_l2075_DUPLICATE_e957_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2069_l2072_l2056_l2075_DUPLICATE_e957_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2056_c2_5cb8_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2056_c2_5cb8_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2056_c2_5cb8_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2056_c2_5cb8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2077_c30_f128_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2075_c7_71b6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2056_c2_5cb8] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2075_c7_71b6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2075_c7_71b6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2075_c7_71b6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2056_c2_5cb8] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2056_c2_5cb8] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output;

     -- t8_MUX[uxn_opcodes_h_l2072_c7_d6ad] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond <= VAR_t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond;
     t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue;
     t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output := t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2056_c2_5cb8] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output;

     -- n8_MUX[uxn_opcodes_h_l2075_c7_71b6] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2075_c7_71b6_cond <= VAR_n8_MUX_uxn_opcodes_h_l2075_c7_71b6_cond;
     n8_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue;
     n8_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output := n8_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output;

     -- MUX[uxn_opcodes_h_l2080_c21_ce84] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l2080_c21_ce84_cond <= VAR_MUX_uxn_opcodes_h_l2080_c21_ce84_cond;
     MUX_uxn_opcodes_h_l2080_c21_ce84_iftrue <= VAR_MUX_uxn_opcodes_h_l2080_c21_ce84_iftrue;
     MUX_uxn_opcodes_h_l2080_c21_ce84_iffalse <= VAR_MUX_uxn_opcodes_h_l2080_c21_ce84_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l2080_c21_ce84_return_output := MUX_uxn_opcodes_h_l2080_c21_ce84_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue := VAR_MUX_uxn_opcodes_h_l2080_c21_ce84_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2072_c7_d6ad] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2072_c7_d6ad] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output;

     -- t8_MUX[uxn_opcodes_h_l2069_c7_fea5] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2069_c7_fea5_cond <= VAR_t8_MUX_uxn_opcodes_h_l2069_c7_fea5_cond;
     t8_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue;
     t8_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output := t8_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output;

     -- n8_MUX[uxn_opcodes_h_l2072_c7_d6ad] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond <= VAR_n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond;
     n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue;
     n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output := n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2075_c7_71b6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output := result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2072_c7_d6ad] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2072_c7_d6ad] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2075_c7_71b6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2069_c7_fea5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2069_c7_fea5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2069_c7_fea5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output;

     -- t8_MUX[uxn_opcodes_h_l2056_c2_5cb8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond <= VAR_t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond;
     t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue;
     t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output := t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2069_c7_fea5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2072_c7_d6ad] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output := result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output;

     -- n8_MUX[uxn_opcodes_h_l2069_c7_fea5] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2069_c7_fea5_cond <= VAR_n8_MUX_uxn_opcodes_h_l2069_c7_fea5_cond;
     n8_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue;
     n8_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output := n8_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2072_c7_d6ad_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2056_c2_5cb8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2056_c2_5cb8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2069_c7_fea5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output := result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2056_c2_5cb8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output;

     -- n8_MUX[uxn_opcodes_h_l2056_c2_5cb8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond <= VAR_n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond;
     n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue;
     n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output := n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2056_c2_5cb8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_fea5_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2056_c2_5cb8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output := result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2052_l2084_DUPLICATE_574d LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2052_l2084_DUPLICATE_574d_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_04b4(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2056_c2_5cb8_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2052_l2084_DUPLICATE_574d_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2052_l2084_DUPLICATE_574d_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
