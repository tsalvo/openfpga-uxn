-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 57
entity ora_0CLK_edc09f97 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ora_0CLK_edc09f97;
architecture arch of ora_0CLK_edc09f97 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1059_c6_c451]
signal BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1059_c2_4f55]
signal n8_MUX_uxn_opcodes_h_l1059_c2_4f55_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1059_c2_4f55]
signal t8_MUX_uxn_opcodes_h_l1059_c2_4f55_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1059_c2_4f55]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1059_c2_4f55]
signal result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1059_c2_4f55]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1059_c2_4f55]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1059_c2_4f55]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1059_c2_4f55]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1064_c11_f2da]
signal BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1064_c7_69bc]
signal n8_MUX_uxn_opcodes_h_l1064_c7_69bc_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1064_c7_69bc]
signal t8_MUX_uxn_opcodes_h_l1064_c7_69bc_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1064_c7_69bc]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1064_c7_69bc]
signal result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1064_c7_69bc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1064_c7_69bc]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1064_c7_69bc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1064_c7_69bc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1067_c11_c029]
signal BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1067_c7_a96b]
signal n8_MUX_uxn_opcodes_h_l1067_c7_a96b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1067_c7_a96b]
signal t8_MUX_uxn_opcodes_h_l1067_c7_a96b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1067_c7_a96b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1067_c7_a96b]
signal result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1067_c7_a96b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1067_c7_a96b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1067_c7_a96b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1067_c7_a96b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1071_c11_51ed]
signal BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1071_c7_571f]
signal n8_MUX_uxn_opcodes_h_l1071_c7_571f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1071_c7_571f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1071_c7_571f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1071_c7_571f]
signal result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1071_c7_571f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1071_c7_571f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1071_c7_571f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1071_c7_571f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1074_c11_2cef]
signal BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1074_c7_1d83]
signal n8_MUX_uxn_opcodes_h_l1074_c7_1d83_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1074_c7_1d83]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1074_c7_1d83]
signal result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1074_c7_1d83]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1074_c7_1d83]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1074_c7_1d83]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1074_c7_1d83]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l1077_c32_5e1a]
signal BIN_OP_AND_uxn_opcodes_h_l1077_c32_5e1a_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1077_c32_5e1a_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1077_c32_5e1a_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1077_c32_c5f5]
signal BIN_OP_GT_uxn_opcodes_h_l1077_c32_c5f5_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1077_c32_c5f5_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1077_c32_c5f5_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1077_c32_5e79]
signal MUX_uxn_opcodes_h_l1077_c32_5e79_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1077_c32_5e79_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1077_c32_5e79_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1077_c32_5e79_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1079_c11_cdd2]
signal BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1079_c7_f1b4]
signal result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1079_c7_f1b4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1079_c7_f1b4]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1079_c7_f1b4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1079_c7_f1b4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output : unsigned(0 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l1083_c24_85d8]
signal BIN_OP_OR_uxn_opcodes_h_l1083_c24_85d8_left : unsigned(7 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l1083_c24_85d8_right : unsigned(7 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l1083_c24_85d8_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1085_c11_317d]
signal BIN_OP_EQ_uxn_opcodes_h_l1085_c11_317d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1085_c11_317d_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1085_c11_317d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1085_c7_899b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1085_c7_899b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_value := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_sp_shift := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.is_opc_done := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451
BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_left,
BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_right,
BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_return_output);

-- n8_MUX_uxn_opcodes_h_l1059_c2_4f55
n8_MUX_uxn_opcodes_h_l1059_c2_4f55 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1059_c2_4f55_cond,
n8_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue,
n8_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse,
n8_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output);

-- t8_MUX_uxn_opcodes_h_l1059_c2_4f55
t8_MUX_uxn_opcodes_h_l1059_c2_4f55 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1059_c2_4f55_cond,
t8_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue,
t8_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse,
t8_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55
result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55
result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_cond,
result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55
result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55
result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55
result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da
BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_left,
BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_right,
BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_return_output);

-- n8_MUX_uxn_opcodes_h_l1064_c7_69bc
n8_MUX_uxn_opcodes_h_l1064_c7_69bc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1064_c7_69bc_cond,
n8_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue,
n8_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse,
n8_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output);

-- t8_MUX_uxn_opcodes_h_l1064_c7_69bc
t8_MUX_uxn_opcodes_h_l1064_c7_69bc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1064_c7_69bc_cond,
t8_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue,
t8_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse,
t8_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc
result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc
result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_cond,
result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc
result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc
result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc
result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029
BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_left,
BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_right,
BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_return_output);

-- n8_MUX_uxn_opcodes_h_l1067_c7_a96b
n8_MUX_uxn_opcodes_h_l1067_c7_a96b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1067_c7_a96b_cond,
n8_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue,
n8_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse,
n8_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output);

-- t8_MUX_uxn_opcodes_h_l1067_c7_a96b
t8_MUX_uxn_opcodes_h_l1067_c7_a96b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1067_c7_a96b_cond,
t8_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue,
t8_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse,
t8_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b
result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_cond,
result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b
result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b
result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b
result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed
BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_left,
BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_right,
BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_return_output);

-- n8_MUX_uxn_opcodes_h_l1071_c7_571f
n8_MUX_uxn_opcodes_h_l1071_c7_571f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1071_c7_571f_cond,
n8_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue,
n8_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse,
n8_MUX_uxn_opcodes_h_l1071_c7_571f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f
result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_cond,
result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f
result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f
result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f
result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef
BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_left,
BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_right,
BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_return_output);

-- n8_MUX_uxn_opcodes_h_l1074_c7_1d83
n8_MUX_uxn_opcodes_h_l1074_c7_1d83 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1074_c7_1d83_cond,
n8_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue,
n8_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse,
n8_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83
result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83
result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_cond,
result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83
result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83
result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83
result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l1077_c32_5e1a
BIN_OP_AND_uxn_opcodes_h_l1077_c32_5e1a : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l1077_c32_5e1a_left,
BIN_OP_AND_uxn_opcodes_h_l1077_c32_5e1a_right,
BIN_OP_AND_uxn_opcodes_h_l1077_c32_5e1a_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1077_c32_c5f5
BIN_OP_GT_uxn_opcodes_h_l1077_c32_c5f5 : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1077_c32_c5f5_left,
BIN_OP_GT_uxn_opcodes_h_l1077_c32_c5f5_right,
BIN_OP_GT_uxn_opcodes_h_l1077_c32_c5f5_return_output);

-- MUX_uxn_opcodes_h_l1077_c32_5e79
MUX_uxn_opcodes_h_l1077_c32_5e79 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1077_c32_5e79_cond,
MUX_uxn_opcodes_h_l1077_c32_5e79_iftrue,
MUX_uxn_opcodes_h_l1077_c32_5e79_iffalse,
MUX_uxn_opcodes_h_l1077_c32_5e79_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2
BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2_left,
BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2_right,
BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4
result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond,
result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4
result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4
result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4
result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l1083_c24_85d8
BIN_OP_OR_uxn_opcodes_h_l1083_c24_85d8 : entity work.BIN_OP_OR_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l1083_c24_85d8_left,
BIN_OP_OR_uxn_opcodes_h_l1083_c24_85d8_right,
BIN_OP_OR_uxn_opcodes_h_l1083_c24_85d8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1085_c11_317d
BIN_OP_EQ_uxn_opcodes_h_l1085_c11_317d : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1085_c11_317d_left,
BIN_OP_EQ_uxn_opcodes_h_l1085_c11_317d_right,
BIN_OP_EQ_uxn_opcodes_h_l1085_c11_317d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b
result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b
result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_return_output,
 n8_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output,
 t8_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_return_output,
 n8_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output,
 t8_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_return_output,
 n8_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output,
 t8_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_return_output,
 n8_MUX_uxn_opcodes_h_l1071_c7_571f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_return_output,
 n8_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output,
 BIN_OP_AND_uxn_opcodes_h_l1077_c32_5e1a_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1077_c32_c5f5_return_output,
 MUX_uxn_opcodes_h_l1077_c32_5e79_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output,
 BIN_OP_OR_uxn_opcodes_h_l1083_c24_85d8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1085_c11_317d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1059_c2_4f55_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1059_c2_4f55_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1061_c3_f5ca : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1064_c7_69bc_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1064_c7_69bc_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1065_c3_f0b6 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1071_c7_571f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1067_c7_a96b_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1067_c7_a96b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1069_c3_3bd1 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1071_c7_571f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1072_c3_db03 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1074_c7_1d83_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1077_c32_5e79_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1077_c32_5e79_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1077_c32_5e79_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1077_c32_5e1a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1077_c32_5e1a_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1077_c32_5e1a_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1077_c32_c5f5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1077_c32_c5f5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1077_c32_c5f5_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1077_c32_5e79_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1082_c3_dcca : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1083_c24_85d8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1083_c24_85d8_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l1083_c24_85d8_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1085_c11_317d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1085_c11_317d_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1085_c11_317d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1074_l1071_l1067_l1064_l1059_DUPLICATE_ba2d_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1079_l1074_l1071_l1067_l1064_l1059_DUPLICATE_a09b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1079_l1071_l1067_l1064_l1059_DUPLICATE_dac7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1074_l1071_l1067_l1064_l1059_l1085_DUPLICATE_0b91_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1079_l1074_l1071_l1067_l1064_l1085_DUPLICATE_f7f4_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1079_l1074_DUPLICATE_dbf6_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l1055_l1090_DUPLICATE_7ee0_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_GT_uxn_opcodes_h_l1077_c32_c5f5_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1061_c3_f5ca := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1061_c3_f5ca;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1065_c3_f0b6 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1065_c3_f0b6;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1069_c3_3bd1 := resize(to_unsigned(2, 2), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1069_c3_3bd1;
     VAR_MUX_uxn_opcodes_h_l1077_c32_5e79_iffalse := resize(to_signed(-1, 2), 8);
     VAR_MUX_uxn_opcodes_h_l1077_c32_5e79_iftrue := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1085_c11_317d_right := to_unsigned(6, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_right := to_unsigned(4, 3);
     VAR_BIN_OP_AND_uxn_opcodes_h_l1077_c32_5e1a_right := to_unsigned(128, 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1072_c3_db03 := resize(to_unsigned(2, 2), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1072_c3_db03;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2_right := to_unsigned(5, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1082_c3_dcca := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1082_c3_dcca;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_BIN_OP_AND_uxn_opcodes_h_l1077_c32_5e1a_left := VAR_ins;
     VAR_BIN_OP_OR_uxn_opcodes_h_l1083_c24_85d8_left := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1085_c11_317d_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_OR_uxn_opcodes_h_l1083_c24_85d8_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1079_l1071_l1067_l1064_l1059_DUPLICATE_dac7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1079_l1071_l1067_l1064_l1059_DUPLICATE_dac7_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1079_l1074_l1071_l1067_l1064_l1085_DUPLICATE_f7f4 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1079_l1074_l1071_l1067_l1064_l1085_DUPLICATE_f7f4_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1059_c6_c451] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_left;
     BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_return_output := BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1079_l1074_DUPLICATE_dbf6 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1079_l1074_DUPLICATE_dbf6_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1064_c11_f2da] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_left;
     BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_return_output := BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1071_c11_51ed] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_left;
     BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_return_output := BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1074_c11_2cef] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_left;
     BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_return_output := BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1079_l1074_l1071_l1067_l1064_l1059_DUPLICATE_a09b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1079_l1074_l1071_l1067_l1064_l1059_DUPLICATE_a09b_return_output := result.stack_value;

     -- BIN_OP_OR[uxn_opcodes_h_l1083_c24_85d8] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l1083_c24_85d8_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l1083_c24_85d8_left;
     BIN_OP_OR_uxn_opcodes_h_l1083_c24_85d8_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l1083_c24_85d8_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l1083_c24_85d8_return_output := BIN_OP_OR_uxn_opcodes_h_l1083_c24_85d8_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1074_l1071_l1067_l1064_l1059_l1085_DUPLICATE_0b91 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1074_l1071_l1067_l1064_l1059_l1085_DUPLICATE_0b91_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1085_c11_317d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1085_c11_317d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1085_c11_317d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1085_c11_317d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1085_c11_317d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1085_c11_317d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1085_c11_317d_return_output;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1074_l1071_l1067_l1064_l1059_DUPLICATE_ba2d LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1074_l1071_l1067_l1064_l1059_DUPLICATE_ba2d_return_output := result.sp_relative_shift;

     -- BIN_OP_AND[uxn_opcodes_h_l1077_c32_5e1a] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l1077_c32_5e1a_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l1077_c32_5e1a_left;
     BIN_OP_AND_uxn_opcodes_h_l1077_c32_5e1a_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l1077_c32_5e1a_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l1077_c32_5e1a_return_output := BIN_OP_AND_uxn_opcodes_h_l1077_c32_5e1a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1067_c11_c029] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_left;
     BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_return_output := BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1079_c11_cdd2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2_left;
     BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2_return_output := BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2_return_output;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l1077_c32_c5f5_left := VAR_BIN_OP_AND_uxn_opcodes_h_l1077_c32_5e1a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1059_c2_4f55_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1059_c2_4f55_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1059_c6_c451_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1064_c7_69bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1064_c7_69bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1064_c11_f2da_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1067_c7_a96b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1067_c7_a96b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1067_c11_c029_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1071_c7_571f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1071_c11_51ed_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1074_c7_1d83_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1074_c11_2cef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1079_c11_cdd2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1085_c11_317d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1085_c11_317d_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l1083_c24_85d8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1074_l1071_l1067_l1064_l1059_DUPLICATE_ba2d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1074_l1071_l1067_l1064_l1059_DUPLICATE_ba2d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1074_l1071_l1067_l1064_l1059_DUPLICATE_ba2d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1074_l1071_l1067_l1064_l1059_DUPLICATE_ba2d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1074_l1071_l1067_l1064_l1059_DUPLICATE_ba2d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1079_l1074_l1071_l1067_l1064_l1085_DUPLICATE_f7f4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1079_l1074_l1071_l1067_l1064_l1085_DUPLICATE_f7f4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1079_l1074_l1071_l1067_l1064_l1085_DUPLICATE_f7f4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1079_l1074_l1071_l1067_l1064_l1085_DUPLICATE_f7f4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1079_l1074_l1071_l1067_l1064_l1085_DUPLICATE_f7f4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1079_l1074_l1071_l1067_l1064_l1085_DUPLICATE_f7f4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1079_l1071_l1067_l1064_l1059_DUPLICATE_dac7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1079_l1071_l1067_l1064_l1059_DUPLICATE_dac7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1079_l1071_l1067_l1064_l1059_DUPLICATE_dac7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1079_l1071_l1067_l1064_l1059_DUPLICATE_dac7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1079_l1071_l1067_l1064_l1059_DUPLICATE_dac7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1074_l1071_l1067_l1064_l1059_l1085_DUPLICATE_0b91_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1074_l1071_l1067_l1064_l1059_l1085_DUPLICATE_0b91_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1074_l1071_l1067_l1064_l1059_l1085_DUPLICATE_0b91_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1074_l1071_l1067_l1064_l1059_l1085_DUPLICATE_0b91_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1074_l1071_l1067_l1064_l1059_l1085_DUPLICATE_0b91_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1074_l1071_l1067_l1064_l1059_l1085_DUPLICATE_0b91_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1079_l1074_DUPLICATE_dbf6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1079_l1074_DUPLICATE_dbf6_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1079_l1074_l1071_l1067_l1064_l1059_DUPLICATE_a09b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1079_l1074_l1071_l1067_l1064_l1059_DUPLICATE_a09b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1079_l1074_l1071_l1067_l1064_l1059_DUPLICATE_a09b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1079_l1074_l1071_l1067_l1064_l1059_DUPLICATE_a09b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1079_l1074_l1071_l1067_l1064_l1059_DUPLICATE_a09b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1079_l1074_l1071_l1067_l1064_l1059_DUPLICATE_a09b_return_output;
     -- result_stack_value_MUX[uxn_opcodes_h_l1079_c7_f1b4] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output := result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1079_c7_f1b4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1085_c7_899b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l1077_c32_c5f5] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1077_c32_c5f5_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1077_c32_c5f5_left;
     BIN_OP_GT_uxn_opcodes_h_l1077_c32_c5f5_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1077_c32_c5f5_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1077_c32_c5f5_return_output := BIN_OP_GT_uxn_opcodes_h_l1077_c32_c5f5_return_output;

     -- n8_MUX[uxn_opcodes_h_l1074_c7_1d83] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1074_c7_1d83_cond <= VAR_n8_MUX_uxn_opcodes_h_l1074_c7_1d83_cond;
     n8_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue;
     n8_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output := n8_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1085_c7_899b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_return_output;

     -- t8_MUX[uxn_opcodes_h_l1067_c7_a96b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1067_c7_a96b_cond <= VAR_t8_MUX_uxn_opcodes_h_l1067_c7_a96b_cond;
     t8_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue;
     t8_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output := t8_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1079_c7_f1b4] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l1077_c32_5e79_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1077_c32_c5f5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1085_c7_899b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1085_c7_899b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1074_c7_1d83] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output;

     -- MUX[uxn_opcodes_h_l1077_c32_5e79] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1077_c32_5e79_cond <= VAR_MUX_uxn_opcodes_h_l1077_c32_5e79_cond;
     MUX_uxn_opcodes_h_l1077_c32_5e79_iftrue <= VAR_MUX_uxn_opcodes_h_l1077_c32_5e79_iftrue;
     MUX_uxn_opcodes_h_l1077_c32_5e79_iffalse <= VAR_MUX_uxn_opcodes_h_l1077_c32_5e79_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1077_c32_5e79_return_output := MUX_uxn_opcodes_h_l1077_c32_5e79_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1074_c7_1d83] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output := result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output;

     -- t8_MUX[uxn_opcodes_h_l1064_c7_69bc] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1064_c7_69bc_cond <= VAR_t8_MUX_uxn_opcodes_h_l1064_c7_69bc_cond;
     t8_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue;
     t8_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output := t8_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1079_c7_f1b4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1074_c7_1d83] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output;

     -- n8_MUX[uxn_opcodes_h_l1071_c7_571f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1071_c7_571f_cond <= VAR_n8_MUX_uxn_opcodes_h_l1071_c7_571f_cond;
     n8_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue;
     n8_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1071_c7_571f_return_output := n8_MUX_uxn_opcodes_h_l1071_c7_571f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1079_c7_f1b4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue := VAR_MUX_uxn_opcodes_h_l1077_c32_5e79_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1071_c7_571f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1079_c7_f1b4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1074_c7_1d83] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output;

     -- t8_MUX[uxn_opcodes_h_l1059_c2_4f55] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1059_c2_4f55_cond <= VAR_t8_MUX_uxn_opcodes_h_l1059_c2_4f55_cond;
     t8_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue;
     t8_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output := t8_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output;

     -- n8_MUX[uxn_opcodes_h_l1067_c7_a96b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1067_c7_a96b_cond <= VAR_n8_MUX_uxn_opcodes_h_l1067_c7_a96b_cond;
     n8_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue;
     n8_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output := n8_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1071_c7_571f] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_return_output := result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1074_c7_1d83] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1071_c7_571f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1074_c7_1d83] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1071_c7_571f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1071_c7_571f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1074_c7_1d83_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1071_c7_571f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1071_c7_571f_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1067_c7_a96b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1071_c7_571f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1071_c7_571f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_return_output;

     -- n8_MUX[uxn_opcodes_h_l1064_c7_69bc] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1064_c7_69bc_cond <= VAR_n8_MUX_uxn_opcodes_h_l1064_c7_69bc_cond;
     n8_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue;
     n8_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output := n8_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1067_c7_a96b] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output := result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1071_c7_571f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1067_c7_a96b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1071_c7_571f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1071_c7_571f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1071_c7_571f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1064_c7_69bc] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1064_c7_69bc] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output := result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1067_c7_a96b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output;

     -- n8_MUX[uxn_opcodes_h_l1059_c2_4f55] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1059_c2_4f55_cond <= VAR_n8_MUX_uxn_opcodes_h_l1059_c2_4f55_cond;
     n8_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue;
     n8_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output := n8_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1067_c7_a96b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1064_c7_69bc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1067_c7_a96b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1067_c7_a96b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1059_c2_4f55] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1064_c7_69bc] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1064_c7_69bc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1059_c2_4f55] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output := result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1064_c7_69bc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1059_c2_4f55] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output;

     -- Submodule level 7
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1064_c7_69bc_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1059_c2_4f55] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1059_c2_4f55] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1059_c2_4f55] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output;

     -- Submodule level 8
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l1055_l1090_DUPLICATE_7ee0 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l1055_l1090_DUPLICATE_7ee0_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1059_c2_4f55_return_output);

     -- Submodule level 9
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l1055_l1090_DUPLICATE_7ee0_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l1055_l1090_DUPLICATE_7ee0_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
