-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 17
entity device_in_0CLK_50065acf is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 device_address : in unsigned(7 downto 0);
 phase : in unsigned(7 downto 0);
 controller0_buttons : in unsigned(7 downto 0);
 previous_device_ram_read : in unsigned(7 downto 0);
 return_output : out device_in_result_t);
end device_in_0CLK_50065acf;
architecture arch of device_in_0CLK_50065acf is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal device : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : device_in_result_t := (
device_ram_address => to_unsigned(0, 8),
dei_value => to_unsigned(0, 8),
is_dei_done => to_unsigned(0, 1))
;
signal REG_COMB_device : unsigned(7 downto 0);
signal REG_COMB_result : device_in_result_t;

-- Each function instance gets signals
-- BIN_OP_AND[uxn_device_h_l396_c11_26dd]
signal BIN_OP_AND_uxn_device_h_l396_c11_26dd_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_device_h_l396_c11_26dd_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_device_h_l396_c11_26dd_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_device_h_l398_c6_e334]
signal BIN_OP_EQ_uxn_device_h_l398_c6_e334_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_device_h_l398_c6_e334_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_device_h_l398_c6_e334_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_device_h_l398_c1_1854]
signal TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_device_h_l401_c7_c00c]
signal FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_device_h_l398_c2_206e]
signal result_MUX_uxn_device_h_l398_c2_206e_cond : unsigned(0 downto 0);
signal result_MUX_uxn_device_h_l398_c2_206e_iftrue : device_in_result_t;
signal result_MUX_uxn_device_h_l398_c2_206e_iffalse : device_in_result_t;
signal result_MUX_uxn_device_h_l398_c2_206e_return_output : device_in_result_t;

-- system_dei[uxn_device_h_l399_c12_1ce4]
signal system_dei_uxn_device_h_l399_c12_1ce4_CLOCK_ENABLE : unsigned(0 downto 0);
signal system_dei_uxn_device_h_l399_c12_1ce4_device_address : unsigned(7 downto 0);
signal system_dei_uxn_device_h_l399_c12_1ce4_phase : unsigned(7 downto 0);
signal system_dei_uxn_device_h_l399_c12_1ce4_previous_device_ram_read : unsigned(7 downto 0);
signal system_dei_uxn_device_h_l399_c12_1ce4_return_output : device_in_result_t;

-- BIN_OP_EQ[uxn_device_h_l401_c11_7730]
signal BIN_OP_EQ_uxn_device_h_l401_c11_7730_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_device_h_l401_c11_7730_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_device_h_l401_c11_7730_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_device_h_l401_c1_11ab]
signal TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_device_h_l404_c7_aaba]
signal FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_device_h_l401_c7_c00c]
signal result_MUX_uxn_device_h_l401_c7_c00c_cond : unsigned(0 downto 0);
signal result_MUX_uxn_device_h_l401_c7_c00c_iftrue : device_in_result_t;
signal result_MUX_uxn_device_h_l401_c7_c00c_iffalse : device_in_result_t;
signal result_MUX_uxn_device_h_l401_c7_c00c_return_output : device_in_result_t;

-- screen_dei[uxn_device_h_l402_c12_10c4]
signal screen_dei_uxn_device_h_l402_c12_10c4_CLOCK_ENABLE : unsigned(0 downto 0);
signal screen_dei_uxn_device_h_l402_c12_10c4_device_address : unsigned(7 downto 0);
signal screen_dei_uxn_device_h_l402_c12_10c4_phase : unsigned(7 downto 0);
signal screen_dei_uxn_device_h_l402_c12_10c4_previous_device_ram_read : unsigned(7 downto 0);
signal screen_dei_uxn_device_h_l402_c12_10c4_return_output : device_in_result_t;

-- BIN_OP_EQ[uxn_device_h_l404_c11_c8ab]
signal BIN_OP_EQ_uxn_device_h_l404_c11_c8ab_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_device_h_l404_c11_c8ab_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_device_h_l404_c11_c8ab_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_device_h_l404_c1_8849]
signal TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_device_h_l407_c1_311f]
signal FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_device_h_l404_c7_aaba]
signal result_MUX_uxn_device_h_l404_c7_aaba_cond : unsigned(0 downto 0);
signal result_MUX_uxn_device_h_l404_c7_aaba_iftrue : device_in_result_t;
signal result_MUX_uxn_device_h_l404_c7_aaba_iffalse : device_in_result_t;
signal result_MUX_uxn_device_h_l404_c7_aaba_return_output : device_in_result_t;

-- controller_dei[uxn_device_h_l405_c12_9489]
signal controller_dei_uxn_device_h_l405_c12_9489_CLOCK_ENABLE : unsigned(0 downto 0);
signal controller_dei_uxn_device_h_l405_c12_9489_device_address : unsigned(7 downto 0);
signal controller_dei_uxn_device_h_l405_c12_9489_phase : unsigned(7 downto 0);
signal controller_dei_uxn_device_h_l405_c12_9489_controller0_buttons : unsigned(7 downto 0);
signal controller_dei_uxn_device_h_l405_c12_9489_previous_device_ram_read : unsigned(7 downto 0);
signal controller_dei_uxn_device_h_l405_c12_9489_return_output : device_in_result_t;

-- generic_dei[uxn_device_h_l408_c12_bddc]
signal generic_dei_uxn_device_h_l408_c12_bddc_CLOCK_ENABLE : unsigned(0 downto 0);
signal generic_dei_uxn_device_h_l408_c12_bddc_device_address : unsigned(7 downto 0);
signal generic_dei_uxn_device_h_l408_c12_bddc_phase : unsigned(7 downto 0);
signal generic_dei_uxn_device_h_l408_c12_bddc_previous_device_ram_read : unsigned(7 downto 0);
signal generic_dei_uxn_device_h_l408_c12_bddc_return_output : device_in_result_t;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_AND_uxn_device_h_l396_c11_26dd
BIN_OP_AND_uxn_device_h_l396_c11_26dd : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_device_h_l396_c11_26dd_left,
BIN_OP_AND_uxn_device_h_l396_c11_26dd_right,
BIN_OP_AND_uxn_device_h_l396_c11_26dd_return_output);

-- BIN_OP_EQ_uxn_device_h_l398_c6_e334
BIN_OP_EQ_uxn_device_h_l398_c6_e334 : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_device_h_l398_c6_e334_left,
BIN_OP_EQ_uxn_device_h_l398_c6_e334_right,
BIN_OP_EQ_uxn_device_h_l398_c6_e334_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854
TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c
FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_return_output);

-- result_MUX_uxn_device_h_l398_c2_206e
result_MUX_uxn_device_h_l398_c2_206e : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
result_MUX_uxn_device_h_l398_c2_206e_cond,
result_MUX_uxn_device_h_l398_c2_206e_iftrue,
result_MUX_uxn_device_h_l398_c2_206e_iffalse,
result_MUX_uxn_device_h_l398_c2_206e_return_output);

-- system_dei_uxn_device_h_l399_c12_1ce4
system_dei_uxn_device_h_l399_c12_1ce4 : entity work.system_dei_0CLK_5e0132c5 port map (
clk,
system_dei_uxn_device_h_l399_c12_1ce4_CLOCK_ENABLE,
system_dei_uxn_device_h_l399_c12_1ce4_device_address,
system_dei_uxn_device_h_l399_c12_1ce4_phase,
system_dei_uxn_device_h_l399_c12_1ce4_previous_device_ram_read,
system_dei_uxn_device_h_l399_c12_1ce4_return_output);

-- BIN_OP_EQ_uxn_device_h_l401_c11_7730
BIN_OP_EQ_uxn_device_h_l401_c11_7730 : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_device_h_l401_c11_7730_left,
BIN_OP_EQ_uxn_device_h_l401_c11_7730_right,
BIN_OP_EQ_uxn_device_h_l401_c11_7730_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab
TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba
FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_return_output);

-- result_MUX_uxn_device_h_l401_c7_c00c
result_MUX_uxn_device_h_l401_c7_c00c : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
result_MUX_uxn_device_h_l401_c7_c00c_cond,
result_MUX_uxn_device_h_l401_c7_c00c_iftrue,
result_MUX_uxn_device_h_l401_c7_c00c_iffalse,
result_MUX_uxn_device_h_l401_c7_c00c_return_output);

-- screen_dei_uxn_device_h_l402_c12_10c4
screen_dei_uxn_device_h_l402_c12_10c4 : entity work.screen_dei_0CLK_d7085478 port map (
clk,
screen_dei_uxn_device_h_l402_c12_10c4_CLOCK_ENABLE,
screen_dei_uxn_device_h_l402_c12_10c4_device_address,
screen_dei_uxn_device_h_l402_c12_10c4_phase,
screen_dei_uxn_device_h_l402_c12_10c4_previous_device_ram_read,
screen_dei_uxn_device_h_l402_c12_10c4_return_output);

-- BIN_OP_EQ_uxn_device_h_l404_c11_c8ab
BIN_OP_EQ_uxn_device_h_l404_c11_c8ab : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_device_h_l404_c11_c8ab_left,
BIN_OP_EQ_uxn_device_h_l404_c11_c8ab_right,
BIN_OP_EQ_uxn_device_h_l404_c11_c8ab_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849
TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f
FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_return_output);

-- result_MUX_uxn_device_h_l404_c7_aaba
result_MUX_uxn_device_h_l404_c7_aaba : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
result_MUX_uxn_device_h_l404_c7_aaba_cond,
result_MUX_uxn_device_h_l404_c7_aaba_iftrue,
result_MUX_uxn_device_h_l404_c7_aaba_iffalse,
result_MUX_uxn_device_h_l404_c7_aaba_return_output);

-- controller_dei_uxn_device_h_l405_c12_9489
controller_dei_uxn_device_h_l405_c12_9489 : entity work.controller_dei_0CLK_b6e68f82 port map (
clk,
controller_dei_uxn_device_h_l405_c12_9489_CLOCK_ENABLE,
controller_dei_uxn_device_h_l405_c12_9489_device_address,
controller_dei_uxn_device_h_l405_c12_9489_phase,
controller_dei_uxn_device_h_l405_c12_9489_controller0_buttons,
controller_dei_uxn_device_h_l405_c12_9489_previous_device_ram_read,
controller_dei_uxn_device_h_l405_c12_9489_return_output);

-- generic_dei_uxn_device_h_l408_c12_bddc
generic_dei_uxn_device_h_l408_c12_bddc : entity work.generic_dei_0CLK_25f4cd11 port map (
clk,
generic_dei_uxn_device_h_l408_c12_bddc_CLOCK_ENABLE,
generic_dei_uxn_device_h_l408_c12_bddc_device_address,
generic_dei_uxn_device_h_l408_c12_bddc_phase,
generic_dei_uxn_device_h_l408_c12_bddc_previous_device_ram_read,
generic_dei_uxn_device_h_l408_c12_bddc_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 device_address,
 phase,
 controller0_buttons,
 previous_device_ram_read,
 -- Registers
 device,
 result,
 -- All submodule outputs
 BIN_OP_AND_uxn_device_h_l396_c11_26dd_return_output,
 BIN_OP_EQ_uxn_device_h_l398_c6_e334_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_return_output,
 result_MUX_uxn_device_h_l398_c2_206e_return_output,
 system_dei_uxn_device_h_l399_c12_1ce4_return_output,
 BIN_OP_EQ_uxn_device_h_l401_c11_7730_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_return_output,
 result_MUX_uxn_device_h_l401_c7_c00c_return_output,
 screen_dei_uxn_device_h_l402_c12_10c4_return_output,
 BIN_OP_EQ_uxn_device_h_l404_c11_c8ab_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_return_output,
 result_MUX_uxn_device_h_l404_c7_aaba_return_output,
 controller_dei_uxn_device_h_l405_c12_9489_return_output,
 generic_dei_uxn_device_h_l408_c12_bddc_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : device_in_result_t;
 variable VAR_device_address : unsigned(7 downto 0);
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_controller0_buttons : unsigned(7 downto 0);
 variable VAR_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_device_h_l396_c11_26dd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_device_h_l396_c11_26dd_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_device_h_l396_c11_26dd_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_device_h_l398_c6_e334_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_device_h_l398_c6_e334_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_device_h_l398_c6_e334_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_device_h_l398_c2_206e_iftrue : device_in_result_t;
 variable VAR_result_MUX_uxn_device_h_l398_c2_206e_iffalse : device_in_result_t;
 variable VAR_result_MUX_uxn_device_h_l401_c7_c00c_return_output : device_in_result_t;
 variable VAR_result_MUX_uxn_device_h_l398_c2_206e_return_output : device_in_result_t;
 variable VAR_result_MUX_uxn_device_h_l398_c2_206e_cond : unsigned(0 downto 0);
 variable VAR_system_dei_uxn_device_h_l399_c12_1ce4_device_address : unsigned(7 downto 0);
 variable VAR_system_dei_uxn_device_h_l399_c12_1ce4_phase : unsigned(7 downto 0);
 variable VAR_system_dei_uxn_device_h_l399_c12_1ce4_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_system_dei_uxn_device_h_l399_c12_1ce4_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_system_dei_uxn_device_h_l399_c12_1ce4_return_output : device_in_result_t;
 variable VAR_BIN_OP_EQ_uxn_device_h_l401_c11_7730_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_device_h_l401_c11_7730_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_device_h_l401_c11_7730_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_device_h_l401_c7_c00c_iftrue : device_in_result_t;
 variable VAR_result_MUX_uxn_device_h_l401_c7_c00c_iffalse : device_in_result_t;
 variable VAR_result_MUX_uxn_device_h_l404_c7_aaba_return_output : device_in_result_t;
 variable VAR_result_MUX_uxn_device_h_l401_c7_c00c_cond : unsigned(0 downto 0);
 variable VAR_screen_dei_uxn_device_h_l402_c12_10c4_device_address : unsigned(7 downto 0);
 variable VAR_screen_dei_uxn_device_h_l402_c12_10c4_phase : unsigned(7 downto 0);
 variable VAR_screen_dei_uxn_device_h_l402_c12_10c4_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_screen_dei_uxn_device_h_l402_c12_10c4_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_screen_dei_uxn_device_h_l402_c12_10c4_return_output : device_in_result_t;
 variable VAR_BIN_OP_EQ_uxn_device_h_l404_c11_c8ab_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_device_h_l404_c11_c8ab_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_device_h_l404_c11_c8ab_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_device_h_l404_c7_aaba_iftrue : device_in_result_t;
 variable VAR_result_MUX_uxn_device_h_l404_c7_aaba_iffalse : device_in_result_t;
 variable VAR_result_MUX_uxn_device_h_l404_c7_aaba_cond : unsigned(0 downto 0);
 variable VAR_controller_dei_uxn_device_h_l405_c12_9489_device_address : unsigned(7 downto 0);
 variable VAR_controller_dei_uxn_device_h_l405_c12_9489_phase : unsigned(7 downto 0);
 variable VAR_controller_dei_uxn_device_h_l405_c12_9489_controller0_buttons : unsigned(7 downto 0);
 variable VAR_controller_dei_uxn_device_h_l405_c12_9489_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_controller_dei_uxn_device_h_l405_c12_9489_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_controller_dei_uxn_device_h_l405_c12_9489_return_output : device_in_result_t;
 variable VAR_generic_dei_uxn_device_h_l408_c12_bddc_device_address : unsigned(7 downto 0);
 variable VAR_generic_dei_uxn_device_h_l408_c12_bddc_phase : unsigned(7 downto 0);
 variable VAR_generic_dei_uxn_device_h_l408_c12_bddc_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_generic_dei_uxn_device_h_l408_c12_bddc_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_generic_dei_uxn_device_h_l408_c12_bddc_return_output : device_in_result_t;
 -- State registers comb logic variables
variable REG_VAR_device : unsigned(7 downto 0);
variable REG_VAR_result : device_in_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_device := device;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_device_h_l404_c11_c8ab_right := to_unsigned(128, 8);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_AND_uxn_device_h_l396_c11_26dd_right := to_unsigned(240, 8);
     VAR_BIN_OP_EQ_uxn_device_h_l401_c11_7730_right := to_unsigned(32, 8);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_device_h_l398_c6_e334_right := to_unsigned(0, 8);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_device_address := device_address;
     VAR_phase := phase;
     VAR_controller0_buttons := controller0_buttons;
     VAR_previous_device_ram_read := previous_device_ram_read;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_iffalse := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_iftrue := VAR_CLOCK_ENABLE;
     VAR_controller_dei_uxn_device_h_l405_c12_9489_controller0_buttons := VAR_controller0_buttons;
     VAR_BIN_OP_AND_uxn_device_h_l396_c11_26dd_left := VAR_device_address;
     VAR_controller_dei_uxn_device_h_l405_c12_9489_device_address := VAR_device_address;
     VAR_generic_dei_uxn_device_h_l408_c12_bddc_device_address := VAR_device_address;
     VAR_screen_dei_uxn_device_h_l402_c12_10c4_device_address := VAR_device_address;
     VAR_system_dei_uxn_device_h_l399_c12_1ce4_device_address := VAR_device_address;
     VAR_controller_dei_uxn_device_h_l405_c12_9489_phase := VAR_phase;
     VAR_generic_dei_uxn_device_h_l408_c12_bddc_phase := VAR_phase;
     VAR_screen_dei_uxn_device_h_l402_c12_10c4_phase := VAR_phase;
     VAR_system_dei_uxn_device_h_l399_c12_1ce4_phase := VAR_phase;
     VAR_controller_dei_uxn_device_h_l405_c12_9489_previous_device_ram_read := VAR_previous_device_ram_read;
     VAR_generic_dei_uxn_device_h_l408_c12_bddc_previous_device_ram_read := VAR_previous_device_ram_read;
     VAR_screen_dei_uxn_device_h_l402_c12_10c4_previous_device_ram_read := VAR_previous_device_ram_read;
     VAR_system_dei_uxn_device_h_l399_c12_1ce4_previous_device_ram_read := VAR_previous_device_ram_read;
     -- BIN_OP_AND[uxn_device_h_l396_c11_26dd] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_device_h_l396_c11_26dd_left <= VAR_BIN_OP_AND_uxn_device_h_l396_c11_26dd_left;
     BIN_OP_AND_uxn_device_h_l396_c11_26dd_right <= VAR_BIN_OP_AND_uxn_device_h_l396_c11_26dd_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_device_h_l396_c11_26dd_return_output := BIN_OP_AND_uxn_device_h_l396_c11_26dd_return_output;

     -- Submodule level 1
     VAR_BIN_OP_EQ_uxn_device_h_l398_c6_e334_left := VAR_BIN_OP_AND_uxn_device_h_l396_c11_26dd_return_output;
     VAR_BIN_OP_EQ_uxn_device_h_l401_c11_7730_left := VAR_BIN_OP_AND_uxn_device_h_l396_c11_26dd_return_output;
     VAR_BIN_OP_EQ_uxn_device_h_l404_c11_c8ab_left := VAR_BIN_OP_AND_uxn_device_h_l396_c11_26dd_return_output;
     REG_VAR_device := VAR_BIN_OP_AND_uxn_device_h_l396_c11_26dd_return_output;
     -- BIN_OP_EQ[uxn_device_h_l398_c6_e334] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_device_h_l398_c6_e334_left <= VAR_BIN_OP_EQ_uxn_device_h_l398_c6_e334_left;
     BIN_OP_EQ_uxn_device_h_l398_c6_e334_right <= VAR_BIN_OP_EQ_uxn_device_h_l398_c6_e334_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_device_h_l398_c6_e334_return_output := BIN_OP_EQ_uxn_device_h_l398_c6_e334_return_output;

     -- BIN_OP_EQ[uxn_device_h_l401_c11_7730] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_device_h_l401_c11_7730_left <= VAR_BIN_OP_EQ_uxn_device_h_l401_c11_7730_left;
     BIN_OP_EQ_uxn_device_h_l401_c11_7730_right <= VAR_BIN_OP_EQ_uxn_device_h_l401_c11_7730_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_device_h_l401_c11_7730_return_output := BIN_OP_EQ_uxn_device_h_l401_c11_7730_return_output;

     -- BIN_OP_EQ[uxn_device_h_l404_c11_c8ab] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_device_h_l404_c11_c8ab_left <= VAR_BIN_OP_EQ_uxn_device_h_l404_c11_c8ab_left;
     BIN_OP_EQ_uxn_device_h_l404_c11_c8ab_right <= VAR_BIN_OP_EQ_uxn_device_h_l404_c11_c8ab_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_device_h_l404_c11_c8ab_return_output := BIN_OP_EQ_uxn_device_h_l404_c11_c8ab_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_cond := VAR_BIN_OP_EQ_uxn_device_h_l398_c6_e334_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_cond := VAR_BIN_OP_EQ_uxn_device_h_l398_c6_e334_return_output;
     VAR_result_MUX_uxn_device_h_l398_c2_206e_cond := VAR_BIN_OP_EQ_uxn_device_h_l398_c6_e334_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_cond := VAR_BIN_OP_EQ_uxn_device_h_l401_c11_7730_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_cond := VAR_BIN_OP_EQ_uxn_device_h_l401_c11_7730_return_output;
     VAR_result_MUX_uxn_device_h_l401_c7_c00c_cond := VAR_BIN_OP_EQ_uxn_device_h_l401_c11_7730_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_cond := VAR_BIN_OP_EQ_uxn_device_h_l404_c11_c8ab_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_cond := VAR_BIN_OP_EQ_uxn_device_h_l404_c11_c8ab_return_output;
     VAR_result_MUX_uxn_device_h_l404_c7_aaba_cond := VAR_BIN_OP_EQ_uxn_device_h_l404_c11_c8ab_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_device_h_l398_c1_1854] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_device_h_l401_c7_c00c] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_return_output;

     -- Submodule level 3
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c7_c00c_return_output;
     VAR_system_dei_uxn_device_h_l399_c12_1ce4_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l398_c1_1854_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_device_h_l404_c7_aaba] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_return_output;

     -- system_dei[uxn_device_h_l399_c12_1ce4] LATENCY=0
     -- Clock enable
     system_dei_uxn_device_h_l399_c12_1ce4_CLOCK_ENABLE <= VAR_system_dei_uxn_device_h_l399_c12_1ce4_CLOCK_ENABLE;
     -- Inputs
     system_dei_uxn_device_h_l399_c12_1ce4_device_address <= VAR_system_dei_uxn_device_h_l399_c12_1ce4_device_address;
     system_dei_uxn_device_h_l399_c12_1ce4_phase <= VAR_system_dei_uxn_device_h_l399_c12_1ce4_phase;
     system_dei_uxn_device_h_l399_c12_1ce4_previous_device_ram_read <= VAR_system_dei_uxn_device_h_l399_c12_1ce4_previous_device_ram_read;
     -- Outputs
     VAR_system_dei_uxn_device_h_l399_c12_1ce4_return_output := system_dei_uxn_device_h_l399_c12_1ce4_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_device_h_l401_c1_11ab] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_return_output;

     -- Submodule level 4
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c7_aaba_return_output;
     VAR_screen_dei_uxn_device_h_l402_c12_10c4_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l401_c1_11ab_return_output;
     VAR_result_MUX_uxn_device_h_l398_c2_206e_iftrue := VAR_system_dei_uxn_device_h_l399_c12_1ce4_return_output;
     -- screen_dei[uxn_device_h_l402_c12_10c4] LATENCY=0
     -- Clock enable
     screen_dei_uxn_device_h_l402_c12_10c4_CLOCK_ENABLE <= VAR_screen_dei_uxn_device_h_l402_c12_10c4_CLOCK_ENABLE;
     -- Inputs
     screen_dei_uxn_device_h_l402_c12_10c4_device_address <= VAR_screen_dei_uxn_device_h_l402_c12_10c4_device_address;
     screen_dei_uxn_device_h_l402_c12_10c4_phase <= VAR_screen_dei_uxn_device_h_l402_c12_10c4_phase;
     screen_dei_uxn_device_h_l402_c12_10c4_previous_device_ram_read <= VAR_screen_dei_uxn_device_h_l402_c12_10c4_previous_device_ram_read;
     -- Outputs
     VAR_screen_dei_uxn_device_h_l402_c12_10c4_return_output := screen_dei_uxn_device_h_l402_c12_10c4_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_device_h_l404_c1_8849] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_device_h_l407_c1_311f] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_return_output;

     -- Submodule level 5
     VAR_generic_dei_uxn_device_h_l408_c12_bddc_CLOCK_ENABLE := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_device_h_l407_c1_311f_return_output;
     VAR_controller_dei_uxn_device_h_l405_c12_9489_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_device_h_l404_c1_8849_return_output;
     VAR_result_MUX_uxn_device_h_l401_c7_c00c_iftrue := VAR_screen_dei_uxn_device_h_l402_c12_10c4_return_output;
     -- controller_dei[uxn_device_h_l405_c12_9489] LATENCY=0
     -- Clock enable
     controller_dei_uxn_device_h_l405_c12_9489_CLOCK_ENABLE <= VAR_controller_dei_uxn_device_h_l405_c12_9489_CLOCK_ENABLE;
     -- Inputs
     controller_dei_uxn_device_h_l405_c12_9489_device_address <= VAR_controller_dei_uxn_device_h_l405_c12_9489_device_address;
     controller_dei_uxn_device_h_l405_c12_9489_phase <= VAR_controller_dei_uxn_device_h_l405_c12_9489_phase;
     controller_dei_uxn_device_h_l405_c12_9489_controller0_buttons <= VAR_controller_dei_uxn_device_h_l405_c12_9489_controller0_buttons;
     controller_dei_uxn_device_h_l405_c12_9489_previous_device_ram_read <= VAR_controller_dei_uxn_device_h_l405_c12_9489_previous_device_ram_read;
     -- Outputs
     VAR_controller_dei_uxn_device_h_l405_c12_9489_return_output := controller_dei_uxn_device_h_l405_c12_9489_return_output;

     -- generic_dei[uxn_device_h_l408_c12_bddc] LATENCY=0
     -- Clock enable
     generic_dei_uxn_device_h_l408_c12_bddc_CLOCK_ENABLE <= VAR_generic_dei_uxn_device_h_l408_c12_bddc_CLOCK_ENABLE;
     -- Inputs
     generic_dei_uxn_device_h_l408_c12_bddc_device_address <= VAR_generic_dei_uxn_device_h_l408_c12_bddc_device_address;
     generic_dei_uxn_device_h_l408_c12_bddc_phase <= VAR_generic_dei_uxn_device_h_l408_c12_bddc_phase;
     generic_dei_uxn_device_h_l408_c12_bddc_previous_device_ram_read <= VAR_generic_dei_uxn_device_h_l408_c12_bddc_previous_device_ram_read;
     -- Outputs
     VAR_generic_dei_uxn_device_h_l408_c12_bddc_return_output := generic_dei_uxn_device_h_l408_c12_bddc_return_output;

     -- Submodule level 6
     VAR_result_MUX_uxn_device_h_l404_c7_aaba_iftrue := VAR_controller_dei_uxn_device_h_l405_c12_9489_return_output;
     VAR_result_MUX_uxn_device_h_l404_c7_aaba_iffalse := VAR_generic_dei_uxn_device_h_l408_c12_bddc_return_output;
     -- result_MUX[uxn_device_h_l404_c7_aaba] LATENCY=0
     -- Inputs
     result_MUX_uxn_device_h_l404_c7_aaba_cond <= VAR_result_MUX_uxn_device_h_l404_c7_aaba_cond;
     result_MUX_uxn_device_h_l404_c7_aaba_iftrue <= VAR_result_MUX_uxn_device_h_l404_c7_aaba_iftrue;
     result_MUX_uxn_device_h_l404_c7_aaba_iffalse <= VAR_result_MUX_uxn_device_h_l404_c7_aaba_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_device_h_l404_c7_aaba_return_output := result_MUX_uxn_device_h_l404_c7_aaba_return_output;

     -- Submodule level 7
     VAR_result_MUX_uxn_device_h_l401_c7_c00c_iffalse := VAR_result_MUX_uxn_device_h_l404_c7_aaba_return_output;
     -- result_MUX[uxn_device_h_l401_c7_c00c] LATENCY=0
     -- Inputs
     result_MUX_uxn_device_h_l401_c7_c00c_cond <= VAR_result_MUX_uxn_device_h_l401_c7_c00c_cond;
     result_MUX_uxn_device_h_l401_c7_c00c_iftrue <= VAR_result_MUX_uxn_device_h_l401_c7_c00c_iftrue;
     result_MUX_uxn_device_h_l401_c7_c00c_iffalse <= VAR_result_MUX_uxn_device_h_l401_c7_c00c_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_device_h_l401_c7_c00c_return_output := result_MUX_uxn_device_h_l401_c7_c00c_return_output;

     -- Submodule level 8
     VAR_result_MUX_uxn_device_h_l398_c2_206e_iffalse := VAR_result_MUX_uxn_device_h_l401_c7_c00c_return_output;
     -- result_MUX[uxn_device_h_l398_c2_206e] LATENCY=0
     -- Inputs
     result_MUX_uxn_device_h_l398_c2_206e_cond <= VAR_result_MUX_uxn_device_h_l398_c2_206e_cond;
     result_MUX_uxn_device_h_l398_c2_206e_iftrue <= VAR_result_MUX_uxn_device_h_l398_c2_206e_iftrue;
     result_MUX_uxn_device_h_l398_c2_206e_iffalse <= VAR_result_MUX_uxn_device_h_l398_c2_206e_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_device_h_l398_c2_206e_return_output := result_MUX_uxn_device_h_l398_c2_206e_return_output;

     -- Submodule level 9
     REG_VAR_result := VAR_result_MUX_uxn_device_h_l398_c2_206e_return_output;
     VAR_return_output := VAR_result_MUX_uxn_device_h_l398_c2_206e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_device <= REG_VAR_device;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     device <= REG_COMB_device;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
