-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 134
entity uint8_mux128_0CLK_9347d63d is
port(
 sel : in unsigned(6 downto 0);
 in0 : in unsigned(7 downto 0);
 in1 : in unsigned(7 downto 0);
 in2 : in unsigned(7 downto 0);
 in3 : in unsigned(7 downto 0);
 in4 : in unsigned(7 downto 0);
 in5 : in unsigned(7 downto 0);
 in6 : in unsigned(7 downto 0);
 in7 : in unsigned(7 downto 0);
 in8 : in unsigned(7 downto 0);
 in9 : in unsigned(7 downto 0);
 in10 : in unsigned(7 downto 0);
 in11 : in unsigned(7 downto 0);
 in12 : in unsigned(7 downto 0);
 in13 : in unsigned(7 downto 0);
 in14 : in unsigned(7 downto 0);
 in15 : in unsigned(7 downto 0);
 in16 : in unsigned(7 downto 0);
 in17 : in unsigned(7 downto 0);
 in18 : in unsigned(7 downto 0);
 in19 : in unsigned(7 downto 0);
 in20 : in unsigned(7 downto 0);
 in21 : in unsigned(7 downto 0);
 in22 : in unsigned(7 downto 0);
 in23 : in unsigned(7 downto 0);
 in24 : in unsigned(7 downto 0);
 in25 : in unsigned(7 downto 0);
 in26 : in unsigned(7 downto 0);
 in27 : in unsigned(7 downto 0);
 in28 : in unsigned(7 downto 0);
 in29 : in unsigned(7 downto 0);
 in30 : in unsigned(7 downto 0);
 in31 : in unsigned(7 downto 0);
 in32 : in unsigned(7 downto 0);
 in33 : in unsigned(7 downto 0);
 in34 : in unsigned(7 downto 0);
 in35 : in unsigned(7 downto 0);
 in36 : in unsigned(7 downto 0);
 in37 : in unsigned(7 downto 0);
 in38 : in unsigned(7 downto 0);
 in39 : in unsigned(7 downto 0);
 in40 : in unsigned(7 downto 0);
 in41 : in unsigned(7 downto 0);
 in42 : in unsigned(7 downto 0);
 in43 : in unsigned(7 downto 0);
 in44 : in unsigned(7 downto 0);
 in45 : in unsigned(7 downto 0);
 in46 : in unsigned(7 downto 0);
 in47 : in unsigned(7 downto 0);
 in48 : in unsigned(7 downto 0);
 in49 : in unsigned(7 downto 0);
 in50 : in unsigned(7 downto 0);
 in51 : in unsigned(7 downto 0);
 in52 : in unsigned(7 downto 0);
 in53 : in unsigned(7 downto 0);
 in54 : in unsigned(7 downto 0);
 in55 : in unsigned(7 downto 0);
 in56 : in unsigned(7 downto 0);
 in57 : in unsigned(7 downto 0);
 in58 : in unsigned(7 downto 0);
 in59 : in unsigned(7 downto 0);
 in60 : in unsigned(7 downto 0);
 in61 : in unsigned(7 downto 0);
 in62 : in unsigned(7 downto 0);
 in63 : in unsigned(7 downto 0);
 in64 : in unsigned(7 downto 0);
 in65 : in unsigned(7 downto 0);
 in66 : in unsigned(7 downto 0);
 in67 : in unsigned(7 downto 0);
 in68 : in unsigned(7 downto 0);
 in69 : in unsigned(7 downto 0);
 in70 : in unsigned(7 downto 0);
 in71 : in unsigned(7 downto 0);
 in72 : in unsigned(7 downto 0);
 in73 : in unsigned(7 downto 0);
 in74 : in unsigned(7 downto 0);
 in75 : in unsigned(7 downto 0);
 in76 : in unsigned(7 downto 0);
 in77 : in unsigned(7 downto 0);
 in78 : in unsigned(7 downto 0);
 in79 : in unsigned(7 downto 0);
 in80 : in unsigned(7 downto 0);
 in81 : in unsigned(7 downto 0);
 in82 : in unsigned(7 downto 0);
 in83 : in unsigned(7 downto 0);
 in84 : in unsigned(7 downto 0);
 in85 : in unsigned(7 downto 0);
 in86 : in unsigned(7 downto 0);
 in87 : in unsigned(7 downto 0);
 in88 : in unsigned(7 downto 0);
 in89 : in unsigned(7 downto 0);
 in90 : in unsigned(7 downto 0);
 in91 : in unsigned(7 downto 0);
 in92 : in unsigned(7 downto 0);
 in93 : in unsigned(7 downto 0);
 in94 : in unsigned(7 downto 0);
 in95 : in unsigned(7 downto 0);
 in96 : in unsigned(7 downto 0);
 in97 : in unsigned(7 downto 0);
 in98 : in unsigned(7 downto 0);
 in99 : in unsigned(7 downto 0);
 in100 : in unsigned(7 downto 0);
 in101 : in unsigned(7 downto 0);
 in102 : in unsigned(7 downto 0);
 in103 : in unsigned(7 downto 0);
 in104 : in unsigned(7 downto 0);
 in105 : in unsigned(7 downto 0);
 in106 : in unsigned(7 downto 0);
 in107 : in unsigned(7 downto 0);
 in108 : in unsigned(7 downto 0);
 in109 : in unsigned(7 downto 0);
 in110 : in unsigned(7 downto 0);
 in111 : in unsigned(7 downto 0);
 in112 : in unsigned(7 downto 0);
 in113 : in unsigned(7 downto 0);
 in114 : in unsigned(7 downto 0);
 in115 : in unsigned(7 downto 0);
 in116 : in unsigned(7 downto 0);
 in117 : in unsigned(7 downto 0);
 in118 : in unsigned(7 downto 0);
 in119 : in unsigned(7 downto 0);
 in120 : in unsigned(7 downto 0);
 in121 : in unsigned(7 downto 0);
 in122 : in unsigned(7 downto 0);
 in123 : in unsigned(7 downto 0);
 in124 : in unsigned(7 downto 0);
 in125 : in unsigned(7 downto 0);
 in126 : in unsigned(7 downto 0);
 in127 : in unsigned(7 downto 0);
 return_output : out unsigned(7 downto 0));
end uint8_mux128_0CLK_9347d63d;
architecture arch of uint8_mux128_0CLK_9347d63d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- layer0_node0_MUX[bit_math_h_l18_c3_5c06]
signal layer0_node0_MUX_bit_math_h_l18_c3_5c06_cond : unsigned(0 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_5c06_iftrue : unsigned(7 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_5c06_iffalse : unsigned(7 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_5c06_return_output : unsigned(7 downto 0);

-- layer0_node1_MUX[bit_math_h_l29_c3_fa46]
signal layer0_node1_MUX_bit_math_h_l29_c3_fa46_cond : unsigned(0 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_fa46_iftrue : unsigned(7 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_fa46_iffalse : unsigned(7 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_fa46_return_output : unsigned(7 downto 0);

-- layer0_node2_MUX[bit_math_h_l40_c3_f68a]
signal layer0_node2_MUX_bit_math_h_l40_c3_f68a_cond : unsigned(0 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_f68a_iftrue : unsigned(7 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_f68a_iffalse : unsigned(7 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_f68a_return_output : unsigned(7 downto 0);

-- layer0_node3_MUX[bit_math_h_l51_c3_b336]
signal layer0_node3_MUX_bit_math_h_l51_c3_b336_cond : unsigned(0 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_b336_iftrue : unsigned(7 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_b336_iffalse : unsigned(7 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_b336_return_output : unsigned(7 downto 0);

-- layer0_node4_MUX[bit_math_h_l62_c3_07e7]
signal layer0_node4_MUX_bit_math_h_l62_c3_07e7_cond : unsigned(0 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_07e7_iftrue : unsigned(7 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_07e7_iffalse : unsigned(7 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_07e7_return_output : unsigned(7 downto 0);

-- layer0_node5_MUX[bit_math_h_l73_c3_282b]
signal layer0_node5_MUX_bit_math_h_l73_c3_282b_cond : unsigned(0 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_282b_iftrue : unsigned(7 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_282b_iffalse : unsigned(7 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_282b_return_output : unsigned(7 downto 0);

-- layer0_node6_MUX[bit_math_h_l84_c3_62f1]
signal layer0_node6_MUX_bit_math_h_l84_c3_62f1_cond : unsigned(0 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_62f1_iftrue : unsigned(7 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_62f1_iffalse : unsigned(7 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_62f1_return_output : unsigned(7 downto 0);

-- layer0_node7_MUX[bit_math_h_l95_c3_567b]
signal layer0_node7_MUX_bit_math_h_l95_c3_567b_cond : unsigned(0 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_567b_iftrue : unsigned(7 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_567b_iffalse : unsigned(7 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_567b_return_output : unsigned(7 downto 0);

-- layer0_node8_MUX[bit_math_h_l106_c3_47e5]
signal layer0_node8_MUX_bit_math_h_l106_c3_47e5_cond : unsigned(0 downto 0);
signal layer0_node8_MUX_bit_math_h_l106_c3_47e5_iftrue : unsigned(7 downto 0);
signal layer0_node8_MUX_bit_math_h_l106_c3_47e5_iffalse : unsigned(7 downto 0);
signal layer0_node8_MUX_bit_math_h_l106_c3_47e5_return_output : unsigned(7 downto 0);

-- layer0_node9_MUX[bit_math_h_l117_c3_f097]
signal layer0_node9_MUX_bit_math_h_l117_c3_f097_cond : unsigned(0 downto 0);
signal layer0_node9_MUX_bit_math_h_l117_c3_f097_iftrue : unsigned(7 downto 0);
signal layer0_node9_MUX_bit_math_h_l117_c3_f097_iffalse : unsigned(7 downto 0);
signal layer0_node9_MUX_bit_math_h_l117_c3_f097_return_output : unsigned(7 downto 0);

-- layer0_node10_MUX[bit_math_h_l128_c3_0e6c]
signal layer0_node10_MUX_bit_math_h_l128_c3_0e6c_cond : unsigned(0 downto 0);
signal layer0_node10_MUX_bit_math_h_l128_c3_0e6c_iftrue : unsigned(7 downto 0);
signal layer0_node10_MUX_bit_math_h_l128_c3_0e6c_iffalse : unsigned(7 downto 0);
signal layer0_node10_MUX_bit_math_h_l128_c3_0e6c_return_output : unsigned(7 downto 0);

-- layer0_node11_MUX[bit_math_h_l139_c3_3ab9]
signal layer0_node11_MUX_bit_math_h_l139_c3_3ab9_cond : unsigned(0 downto 0);
signal layer0_node11_MUX_bit_math_h_l139_c3_3ab9_iftrue : unsigned(7 downto 0);
signal layer0_node11_MUX_bit_math_h_l139_c3_3ab9_iffalse : unsigned(7 downto 0);
signal layer0_node11_MUX_bit_math_h_l139_c3_3ab9_return_output : unsigned(7 downto 0);

-- layer0_node12_MUX[bit_math_h_l150_c3_e611]
signal layer0_node12_MUX_bit_math_h_l150_c3_e611_cond : unsigned(0 downto 0);
signal layer0_node12_MUX_bit_math_h_l150_c3_e611_iftrue : unsigned(7 downto 0);
signal layer0_node12_MUX_bit_math_h_l150_c3_e611_iffalse : unsigned(7 downto 0);
signal layer0_node12_MUX_bit_math_h_l150_c3_e611_return_output : unsigned(7 downto 0);

-- layer0_node13_MUX[bit_math_h_l161_c3_e037]
signal layer0_node13_MUX_bit_math_h_l161_c3_e037_cond : unsigned(0 downto 0);
signal layer0_node13_MUX_bit_math_h_l161_c3_e037_iftrue : unsigned(7 downto 0);
signal layer0_node13_MUX_bit_math_h_l161_c3_e037_iffalse : unsigned(7 downto 0);
signal layer0_node13_MUX_bit_math_h_l161_c3_e037_return_output : unsigned(7 downto 0);

-- layer0_node14_MUX[bit_math_h_l172_c3_ad25]
signal layer0_node14_MUX_bit_math_h_l172_c3_ad25_cond : unsigned(0 downto 0);
signal layer0_node14_MUX_bit_math_h_l172_c3_ad25_iftrue : unsigned(7 downto 0);
signal layer0_node14_MUX_bit_math_h_l172_c3_ad25_iffalse : unsigned(7 downto 0);
signal layer0_node14_MUX_bit_math_h_l172_c3_ad25_return_output : unsigned(7 downto 0);

-- layer0_node15_MUX[bit_math_h_l183_c3_dacd]
signal layer0_node15_MUX_bit_math_h_l183_c3_dacd_cond : unsigned(0 downto 0);
signal layer0_node15_MUX_bit_math_h_l183_c3_dacd_iftrue : unsigned(7 downto 0);
signal layer0_node15_MUX_bit_math_h_l183_c3_dacd_iffalse : unsigned(7 downto 0);
signal layer0_node15_MUX_bit_math_h_l183_c3_dacd_return_output : unsigned(7 downto 0);

-- layer0_node16_MUX[bit_math_h_l194_c3_5393]
signal layer0_node16_MUX_bit_math_h_l194_c3_5393_cond : unsigned(0 downto 0);
signal layer0_node16_MUX_bit_math_h_l194_c3_5393_iftrue : unsigned(7 downto 0);
signal layer0_node16_MUX_bit_math_h_l194_c3_5393_iffalse : unsigned(7 downto 0);
signal layer0_node16_MUX_bit_math_h_l194_c3_5393_return_output : unsigned(7 downto 0);

-- layer0_node17_MUX[bit_math_h_l205_c3_4246]
signal layer0_node17_MUX_bit_math_h_l205_c3_4246_cond : unsigned(0 downto 0);
signal layer0_node17_MUX_bit_math_h_l205_c3_4246_iftrue : unsigned(7 downto 0);
signal layer0_node17_MUX_bit_math_h_l205_c3_4246_iffalse : unsigned(7 downto 0);
signal layer0_node17_MUX_bit_math_h_l205_c3_4246_return_output : unsigned(7 downto 0);

-- layer0_node18_MUX[bit_math_h_l216_c3_2748]
signal layer0_node18_MUX_bit_math_h_l216_c3_2748_cond : unsigned(0 downto 0);
signal layer0_node18_MUX_bit_math_h_l216_c3_2748_iftrue : unsigned(7 downto 0);
signal layer0_node18_MUX_bit_math_h_l216_c3_2748_iffalse : unsigned(7 downto 0);
signal layer0_node18_MUX_bit_math_h_l216_c3_2748_return_output : unsigned(7 downto 0);

-- layer0_node19_MUX[bit_math_h_l227_c3_1dae]
signal layer0_node19_MUX_bit_math_h_l227_c3_1dae_cond : unsigned(0 downto 0);
signal layer0_node19_MUX_bit_math_h_l227_c3_1dae_iftrue : unsigned(7 downto 0);
signal layer0_node19_MUX_bit_math_h_l227_c3_1dae_iffalse : unsigned(7 downto 0);
signal layer0_node19_MUX_bit_math_h_l227_c3_1dae_return_output : unsigned(7 downto 0);

-- layer0_node20_MUX[bit_math_h_l238_c3_e7c7]
signal layer0_node20_MUX_bit_math_h_l238_c3_e7c7_cond : unsigned(0 downto 0);
signal layer0_node20_MUX_bit_math_h_l238_c3_e7c7_iftrue : unsigned(7 downto 0);
signal layer0_node20_MUX_bit_math_h_l238_c3_e7c7_iffalse : unsigned(7 downto 0);
signal layer0_node20_MUX_bit_math_h_l238_c3_e7c7_return_output : unsigned(7 downto 0);

-- layer0_node21_MUX[bit_math_h_l249_c3_8f8c]
signal layer0_node21_MUX_bit_math_h_l249_c3_8f8c_cond : unsigned(0 downto 0);
signal layer0_node21_MUX_bit_math_h_l249_c3_8f8c_iftrue : unsigned(7 downto 0);
signal layer0_node21_MUX_bit_math_h_l249_c3_8f8c_iffalse : unsigned(7 downto 0);
signal layer0_node21_MUX_bit_math_h_l249_c3_8f8c_return_output : unsigned(7 downto 0);

-- layer0_node22_MUX[bit_math_h_l260_c3_321e]
signal layer0_node22_MUX_bit_math_h_l260_c3_321e_cond : unsigned(0 downto 0);
signal layer0_node22_MUX_bit_math_h_l260_c3_321e_iftrue : unsigned(7 downto 0);
signal layer0_node22_MUX_bit_math_h_l260_c3_321e_iffalse : unsigned(7 downto 0);
signal layer0_node22_MUX_bit_math_h_l260_c3_321e_return_output : unsigned(7 downto 0);

-- layer0_node23_MUX[bit_math_h_l271_c3_86c3]
signal layer0_node23_MUX_bit_math_h_l271_c3_86c3_cond : unsigned(0 downto 0);
signal layer0_node23_MUX_bit_math_h_l271_c3_86c3_iftrue : unsigned(7 downto 0);
signal layer0_node23_MUX_bit_math_h_l271_c3_86c3_iffalse : unsigned(7 downto 0);
signal layer0_node23_MUX_bit_math_h_l271_c3_86c3_return_output : unsigned(7 downto 0);

-- layer0_node24_MUX[bit_math_h_l282_c3_2992]
signal layer0_node24_MUX_bit_math_h_l282_c3_2992_cond : unsigned(0 downto 0);
signal layer0_node24_MUX_bit_math_h_l282_c3_2992_iftrue : unsigned(7 downto 0);
signal layer0_node24_MUX_bit_math_h_l282_c3_2992_iffalse : unsigned(7 downto 0);
signal layer0_node24_MUX_bit_math_h_l282_c3_2992_return_output : unsigned(7 downto 0);

-- layer0_node25_MUX[bit_math_h_l293_c3_ece2]
signal layer0_node25_MUX_bit_math_h_l293_c3_ece2_cond : unsigned(0 downto 0);
signal layer0_node25_MUX_bit_math_h_l293_c3_ece2_iftrue : unsigned(7 downto 0);
signal layer0_node25_MUX_bit_math_h_l293_c3_ece2_iffalse : unsigned(7 downto 0);
signal layer0_node25_MUX_bit_math_h_l293_c3_ece2_return_output : unsigned(7 downto 0);

-- layer0_node26_MUX[bit_math_h_l304_c3_7f9b]
signal layer0_node26_MUX_bit_math_h_l304_c3_7f9b_cond : unsigned(0 downto 0);
signal layer0_node26_MUX_bit_math_h_l304_c3_7f9b_iftrue : unsigned(7 downto 0);
signal layer0_node26_MUX_bit_math_h_l304_c3_7f9b_iffalse : unsigned(7 downto 0);
signal layer0_node26_MUX_bit_math_h_l304_c3_7f9b_return_output : unsigned(7 downto 0);

-- layer0_node27_MUX[bit_math_h_l315_c3_5c0f]
signal layer0_node27_MUX_bit_math_h_l315_c3_5c0f_cond : unsigned(0 downto 0);
signal layer0_node27_MUX_bit_math_h_l315_c3_5c0f_iftrue : unsigned(7 downto 0);
signal layer0_node27_MUX_bit_math_h_l315_c3_5c0f_iffalse : unsigned(7 downto 0);
signal layer0_node27_MUX_bit_math_h_l315_c3_5c0f_return_output : unsigned(7 downto 0);

-- layer0_node28_MUX[bit_math_h_l326_c3_12a3]
signal layer0_node28_MUX_bit_math_h_l326_c3_12a3_cond : unsigned(0 downto 0);
signal layer0_node28_MUX_bit_math_h_l326_c3_12a3_iftrue : unsigned(7 downto 0);
signal layer0_node28_MUX_bit_math_h_l326_c3_12a3_iffalse : unsigned(7 downto 0);
signal layer0_node28_MUX_bit_math_h_l326_c3_12a3_return_output : unsigned(7 downto 0);

-- layer0_node29_MUX[bit_math_h_l337_c3_cbb8]
signal layer0_node29_MUX_bit_math_h_l337_c3_cbb8_cond : unsigned(0 downto 0);
signal layer0_node29_MUX_bit_math_h_l337_c3_cbb8_iftrue : unsigned(7 downto 0);
signal layer0_node29_MUX_bit_math_h_l337_c3_cbb8_iffalse : unsigned(7 downto 0);
signal layer0_node29_MUX_bit_math_h_l337_c3_cbb8_return_output : unsigned(7 downto 0);

-- layer0_node30_MUX[bit_math_h_l348_c3_8c5c]
signal layer0_node30_MUX_bit_math_h_l348_c3_8c5c_cond : unsigned(0 downto 0);
signal layer0_node30_MUX_bit_math_h_l348_c3_8c5c_iftrue : unsigned(7 downto 0);
signal layer0_node30_MUX_bit_math_h_l348_c3_8c5c_iffalse : unsigned(7 downto 0);
signal layer0_node30_MUX_bit_math_h_l348_c3_8c5c_return_output : unsigned(7 downto 0);

-- layer0_node31_MUX[bit_math_h_l359_c3_d6b9]
signal layer0_node31_MUX_bit_math_h_l359_c3_d6b9_cond : unsigned(0 downto 0);
signal layer0_node31_MUX_bit_math_h_l359_c3_d6b9_iftrue : unsigned(7 downto 0);
signal layer0_node31_MUX_bit_math_h_l359_c3_d6b9_iffalse : unsigned(7 downto 0);
signal layer0_node31_MUX_bit_math_h_l359_c3_d6b9_return_output : unsigned(7 downto 0);

-- layer0_node32_MUX[bit_math_h_l370_c3_3d24]
signal layer0_node32_MUX_bit_math_h_l370_c3_3d24_cond : unsigned(0 downto 0);
signal layer0_node32_MUX_bit_math_h_l370_c3_3d24_iftrue : unsigned(7 downto 0);
signal layer0_node32_MUX_bit_math_h_l370_c3_3d24_iffalse : unsigned(7 downto 0);
signal layer0_node32_MUX_bit_math_h_l370_c3_3d24_return_output : unsigned(7 downto 0);

-- layer0_node33_MUX[bit_math_h_l381_c3_bdd0]
signal layer0_node33_MUX_bit_math_h_l381_c3_bdd0_cond : unsigned(0 downto 0);
signal layer0_node33_MUX_bit_math_h_l381_c3_bdd0_iftrue : unsigned(7 downto 0);
signal layer0_node33_MUX_bit_math_h_l381_c3_bdd0_iffalse : unsigned(7 downto 0);
signal layer0_node33_MUX_bit_math_h_l381_c3_bdd0_return_output : unsigned(7 downto 0);

-- layer0_node34_MUX[bit_math_h_l392_c3_f617]
signal layer0_node34_MUX_bit_math_h_l392_c3_f617_cond : unsigned(0 downto 0);
signal layer0_node34_MUX_bit_math_h_l392_c3_f617_iftrue : unsigned(7 downto 0);
signal layer0_node34_MUX_bit_math_h_l392_c3_f617_iffalse : unsigned(7 downto 0);
signal layer0_node34_MUX_bit_math_h_l392_c3_f617_return_output : unsigned(7 downto 0);

-- layer0_node35_MUX[bit_math_h_l403_c3_683e]
signal layer0_node35_MUX_bit_math_h_l403_c3_683e_cond : unsigned(0 downto 0);
signal layer0_node35_MUX_bit_math_h_l403_c3_683e_iftrue : unsigned(7 downto 0);
signal layer0_node35_MUX_bit_math_h_l403_c3_683e_iffalse : unsigned(7 downto 0);
signal layer0_node35_MUX_bit_math_h_l403_c3_683e_return_output : unsigned(7 downto 0);

-- layer0_node36_MUX[bit_math_h_l414_c3_cd2c]
signal layer0_node36_MUX_bit_math_h_l414_c3_cd2c_cond : unsigned(0 downto 0);
signal layer0_node36_MUX_bit_math_h_l414_c3_cd2c_iftrue : unsigned(7 downto 0);
signal layer0_node36_MUX_bit_math_h_l414_c3_cd2c_iffalse : unsigned(7 downto 0);
signal layer0_node36_MUX_bit_math_h_l414_c3_cd2c_return_output : unsigned(7 downto 0);

-- layer0_node37_MUX[bit_math_h_l425_c3_2485]
signal layer0_node37_MUX_bit_math_h_l425_c3_2485_cond : unsigned(0 downto 0);
signal layer0_node37_MUX_bit_math_h_l425_c3_2485_iftrue : unsigned(7 downto 0);
signal layer0_node37_MUX_bit_math_h_l425_c3_2485_iffalse : unsigned(7 downto 0);
signal layer0_node37_MUX_bit_math_h_l425_c3_2485_return_output : unsigned(7 downto 0);

-- layer0_node38_MUX[bit_math_h_l436_c3_c940]
signal layer0_node38_MUX_bit_math_h_l436_c3_c940_cond : unsigned(0 downto 0);
signal layer0_node38_MUX_bit_math_h_l436_c3_c940_iftrue : unsigned(7 downto 0);
signal layer0_node38_MUX_bit_math_h_l436_c3_c940_iffalse : unsigned(7 downto 0);
signal layer0_node38_MUX_bit_math_h_l436_c3_c940_return_output : unsigned(7 downto 0);

-- layer0_node39_MUX[bit_math_h_l447_c3_b150]
signal layer0_node39_MUX_bit_math_h_l447_c3_b150_cond : unsigned(0 downto 0);
signal layer0_node39_MUX_bit_math_h_l447_c3_b150_iftrue : unsigned(7 downto 0);
signal layer0_node39_MUX_bit_math_h_l447_c3_b150_iffalse : unsigned(7 downto 0);
signal layer0_node39_MUX_bit_math_h_l447_c3_b150_return_output : unsigned(7 downto 0);

-- layer0_node40_MUX[bit_math_h_l458_c3_c977]
signal layer0_node40_MUX_bit_math_h_l458_c3_c977_cond : unsigned(0 downto 0);
signal layer0_node40_MUX_bit_math_h_l458_c3_c977_iftrue : unsigned(7 downto 0);
signal layer0_node40_MUX_bit_math_h_l458_c3_c977_iffalse : unsigned(7 downto 0);
signal layer0_node40_MUX_bit_math_h_l458_c3_c977_return_output : unsigned(7 downto 0);

-- layer0_node41_MUX[bit_math_h_l469_c3_b3bf]
signal layer0_node41_MUX_bit_math_h_l469_c3_b3bf_cond : unsigned(0 downto 0);
signal layer0_node41_MUX_bit_math_h_l469_c3_b3bf_iftrue : unsigned(7 downto 0);
signal layer0_node41_MUX_bit_math_h_l469_c3_b3bf_iffalse : unsigned(7 downto 0);
signal layer0_node41_MUX_bit_math_h_l469_c3_b3bf_return_output : unsigned(7 downto 0);

-- layer0_node42_MUX[bit_math_h_l480_c3_c677]
signal layer0_node42_MUX_bit_math_h_l480_c3_c677_cond : unsigned(0 downto 0);
signal layer0_node42_MUX_bit_math_h_l480_c3_c677_iftrue : unsigned(7 downto 0);
signal layer0_node42_MUX_bit_math_h_l480_c3_c677_iffalse : unsigned(7 downto 0);
signal layer0_node42_MUX_bit_math_h_l480_c3_c677_return_output : unsigned(7 downto 0);

-- layer0_node43_MUX[bit_math_h_l491_c3_2838]
signal layer0_node43_MUX_bit_math_h_l491_c3_2838_cond : unsigned(0 downto 0);
signal layer0_node43_MUX_bit_math_h_l491_c3_2838_iftrue : unsigned(7 downto 0);
signal layer0_node43_MUX_bit_math_h_l491_c3_2838_iffalse : unsigned(7 downto 0);
signal layer0_node43_MUX_bit_math_h_l491_c3_2838_return_output : unsigned(7 downto 0);

-- layer0_node44_MUX[bit_math_h_l502_c3_6b96]
signal layer0_node44_MUX_bit_math_h_l502_c3_6b96_cond : unsigned(0 downto 0);
signal layer0_node44_MUX_bit_math_h_l502_c3_6b96_iftrue : unsigned(7 downto 0);
signal layer0_node44_MUX_bit_math_h_l502_c3_6b96_iffalse : unsigned(7 downto 0);
signal layer0_node44_MUX_bit_math_h_l502_c3_6b96_return_output : unsigned(7 downto 0);

-- layer0_node45_MUX[bit_math_h_l513_c3_b86e]
signal layer0_node45_MUX_bit_math_h_l513_c3_b86e_cond : unsigned(0 downto 0);
signal layer0_node45_MUX_bit_math_h_l513_c3_b86e_iftrue : unsigned(7 downto 0);
signal layer0_node45_MUX_bit_math_h_l513_c3_b86e_iffalse : unsigned(7 downto 0);
signal layer0_node45_MUX_bit_math_h_l513_c3_b86e_return_output : unsigned(7 downto 0);

-- layer0_node46_MUX[bit_math_h_l524_c3_4ef5]
signal layer0_node46_MUX_bit_math_h_l524_c3_4ef5_cond : unsigned(0 downto 0);
signal layer0_node46_MUX_bit_math_h_l524_c3_4ef5_iftrue : unsigned(7 downto 0);
signal layer0_node46_MUX_bit_math_h_l524_c3_4ef5_iffalse : unsigned(7 downto 0);
signal layer0_node46_MUX_bit_math_h_l524_c3_4ef5_return_output : unsigned(7 downto 0);

-- layer0_node47_MUX[bit_math_h_l535_c3_21f3]
signal layer0_node47_MUX_bit_math_h_l535_c3_21f3_cond : unsigned(0 downto 0);
signal layer0_node47_MUX_bit_math_h_l535_c3_21f3_iftrue : unsigned(7 downto 0);
signal layer0_node47_MUX_bit_math_h_l535_c3_21f3_iffalse : unsigned(7 downto 0);
signal layer0_node47_MUX_bit_math_h_l535_c3_21f3_return_output : unsigned(7 downto 0);

-- layer0_node48_MUX[bit_math_h_l546_c3_5be4]
signal layer0_node48_MUX_bit_math_h_l546_c3_5be4_cond : unsigned(0 downto 0);
signal layer0_node48_MUX_bit_math_h_l546_c3_5be4_iftrue : unsigned(7 downto 0);
signal layer0_node48_MUX_bit_math_h_l546_c3_5be4_iffalse : unsigned(7 downto 0);
signal layer0_node48_MUX_bit_math_h_l546_c3_5be4_return_output : unsigned(7 downto 0);

-- layer0_node49_MUX[bit_math_h_l557_c3_3410]
signal layer0_node49_MUX_bit_math_h_l557_c3_3410_cond : unsigned(0 downto 0);
signal layer0_node49_MUX_bit_math_h_l557_c3_3410_iftrue : unsigned(7 downto 0);
signal layer0_node49_MUX_bit_math_h_l557_c3_3410_iffalse : unsigned(7 downto 0);
signal layer0_node49_MUX_bit_math_h_l557_c3_3410_return_output : unsigned(7 downto 0);

-- layer0_node50_MUX[bit_math_h_l568_c3_4522]
signal layer0_node50_MUX_bit_math_h_l568_c3_4522_cond : unsigned(0 downto 0);
signal layer0_node50_MUX_bit_math_h_l568_c3_4522_iftrue : unsigned(7 downto 0);
signal layer0_node50_MUX_bit_math_h_l568_c3_4522_iffalse : unsigned(7 downto 0);
signal layer0_node50_MUX_bit_math_h_l568_c3_4522_return_output : unsigned(7 downto 0);

-- layer0_node51_MUX[bit_math_h_l579_c3_8398]
signal layer0_node51_MUX_bit_math_h_l579_c3_8398_cond : unsigned(0 downto 0);
signal layer0_node51_MUX_bit_math_h_l579_c3_8398_iftrue : unsigned(7 downto 0);
signal layer0_node51_MUX_bit_math_h_l579_c3_8398_iffalse : unsigned(7 downto 0);
signal layer0_node51_MUX_bit_math_h_l579_c3_8398_return_output : unsigned(7 downto 0);

-- layer0_node52_MUX[bit_math_h_l590_c3_6d3d]
signal layer0_node52_MUX_bit_math_h_l590_c3_6d3d_cond : unsigned(0 downto 0);
signal layer0_node52_MUX_bit_math_h_l590_c3_6d3d_iftrue : unsigned(7 downto 0);
signal layer0_node52_MUX_bit_math_h_l590_c3_6d3d_iffalse : unsigned(7 downto 0);
signal layer0_node52_MUX_bit_math_h_l590_c3_6d3d_return_output : unsigned(7 downto 0);

-- layer0_node53_MUX[bit_math_h_l601_c3_6dc2]
signal layer0_node53_MUX_bit_math_h_l601_c3_6dc2_cond : unsigned(0 downto 0);
signal layer0_node53_MUX_bit_math_h_l601_c3_6dc2_iftrue : unsigned(7 downto 0);
signal layer0_node53_MUX_bit_math_h_l601_c3_6dc2_iffalse : unsigned(7 downto 0);
signal layer0_node53_MUX_bit_math_h_l601_c3_6dc2_return_output : unsigned(7 downto 0);

-- layer0_node54_MUX[bit_math_h_l612_c3_cab9]
signal layer0_node54_MUX_bit_math_h_l612_c3_cab9_cond : unsigned(0 downto 0);
signal layer0_node54_MUX_bit_math_h_l612_c3_cab9_iftrue : unsigned(7 downto 0);
signal layer0_node54_MUX_bit_math_h_l612_c3_cab9_iffalse : unsigned(7 downto 0);
signal layer0_node54_MUX_bit_math_h_l612_c3_cab9_return_output : unsigned(7 downto 0);

-- layer0_node55_MUX[bit_math_h_l623_c3_2e5e]
signal layer0_node55_MUX_bit_math_h_l623_c3_2e5e_cond : unsigned(0 downto 0);
signal layer0_node55_MUX_bit_math_h_l623_c3_2e5e_iftrue : unsigned(7 downto 0);
signal layer0_node55_MUX_bit_math_h_l623_c3_2e5e_iffalse : unsigned(7 downto 0);
signal layer0_node55_MUX_bit_math_h_l623_c3_2e5e_return_output : unsigned(7 downto 0);

-- layer0_node56_MUX[bit_math_h_l634_c3_ab19]
signal layer0_node56_MUX_bit_math_h_l634_c3_ab19_cond : unsigned(0 downto 0);
signal layer0_node56_MUX_bit_math_h_l634_c3_ab19_iftrue : unsigned(7 downto 0);
signal layer0_node56_MUX_bit_math_h_l634_c3_ab19_iffalse : unsigned(7 downto 0);
signal layer0_node56_MUX_bit_math_h_l634_c3_ab19_return_output : unsigned(7 downto 0);

-- layer0_node57_MUX[bit_math_h_l645_c3_cec5]
signal layer0_node57_MUX_bit_math_h_l645_c3_cec5_cond : unsigned(0 downto 0);
signal layer0_node57_MUX_bit_math_h_l645_c3_cec5_iftrue : unsigned(7 downto 0);
signal layer0_node57_MUX_bit_math_h_l645_c3_cec5_iffalse : unsigned(7 downto 0);
signal layer0_node57_MUX_bit_math_h_l645_c3_cec5_return_output : unsigned(7 downto 0);

-- layer0_node58_MUX[bit_math_h_l656_c3_312b]
signal layer0_node58_MUX_bit_math_h_l656_c3_312b_cond : unsigned(0 downto 0);
signal layer0_node58_MUX_bit_math_h_l656_c3_312b_iftrue : unsigned(7 downto 0);
signal layer0_node58_MUX_bit_math_h_l656_c3_312b_iffalse : unsigned(7 downto 0);
signal layer0_node58_MUX_bit_math_h_l656_c3_312b_return_output : unsigned(7 downto 0);

-- layer0_node59_MUX[bit_math_h_l667_c3_672d]
signal layer0_node59_MUX_bit_math_h_l667_c3_672d_cond : unsigned(0 downto 0);
signal layer0_node59_MUX_bit_math_h_l667_c3_672d_iftrue : unsigned(7 downto 0);
signal layer0_node59_MUX_bit_math_h_l667_c3_672d_iffalse : unsigned(7 downto 0);
signal layer0_node59_MUX_bit_math_h_l667_c3_672d_return_output : unsigned(7 downto 0);

-- layer0_node60_MUX[bit_math_h_l678_c3_9a42]
signal layer0_node60_MUX_bit_math_h_l678_c3_9a42_cond : unsigned(0 downto 0);
signal layer0_node60_MUX_bit_math_h_l678_c3_9a42_iftrue : unsigned(7 downto 0);
signal layer0_node60_MUX_bit_math_h_l678_c3_9a42_iffalse : unsigned(7 downto 0);
signal layer0_node60_MUX_bit_math_h_l678_c3_9a42_return_output : unsigned(7 downto 0);

-- layer0_node61_MUX[bit_math_h_l689_c3_be95]
signal layer0_node61_MUX_bit_math_h_l689_c3_be95_cond : unsigned(0 downto 0);
signal layer0_node61_MUX_bit_math_h_l689_c3_be95_iftrue : unsigned(7 downto 0);
signal layer0_node61_MUX_bit_math_h_l689_c3_be95_iffalse : unsigned(7 downto 0);
signal layer0_node61_MUX_bit_math_h_l689_c3_be95_return_output : unsigned(7 downto 0);

-- layer0_node62_MUX[bit_math_h_l700_c3_8a98]
signal layer0_node62_MUX_bit_math_h_l700_c3_8a98_cond : unsigned(0 downto 0);
signal layer0_node62_MUX_bit_math_h_l700_c3_8a98_iftrue : unsigned(7 downto 0);
signal layer0_node62_MUX_bit_math_h_l700_c3_8a98_iffalse : unsigned(7 downto 0);
signal layer0_node62_MUX_bit_math_h_l700_c3_8a98_return_output : unsigned(7 downto 0);

-- layer0_node63_MUX[bit_math_h_l711_c3_45fc]
signal layer0_node63_MUX_bit_math_h_l711_c3_45fc_cond : unsigned(0 downto 0);
signal layer0_node63_MUX_bit_math_h_l711_c3_45fc_iftrue : unsigned(7 downto 0);
signal layer0_node63_MUX_bit_math_h_l711_c3_45fc_iffalse : unsigned(7 downto 0);
signal layer0_node63_MUX_bit_math_h_l711_c3_45fc_return_output : unsigned(7 downto 0);

-- layer1_node0_MUX[bit_math_h_l728_c3_2ff0]
signal layer1_node0_MUX_bit_math_h_l728_c3_2ff0_cond : unsigned(0 downto 0);
signal layer1_node0_MUX_bit_math_h_l728_c3_2ff0_iftrue : unsigned(7 downto 0);
signal layer1_node0_MUX_bit_math_h_l728_c3_2ff0_iffalse : unsigned(7 downto 0);
signal layer1_node0_MUX_bit_math_h_l728_c3_2ff0_return_output : unsigned(7 downto 0);

-- layer1_node1_MUX[bit_math_h_l739_c3_8d8d]
signal layer1_node1_MUX_bit_math_h_l739_c3_8d8d_cond : unsigned(0 downto 0);
signal layer1_node1_MUX_bit_math_h_l739_c3_8d8d_iftrue : unsigned(7 downto 0);
signal layer1_node1_MUX_bit_math_h_l739_c3_8d8d_iffalse : unsigned(7 downto 0);
signal layer1_node1_MUX_bit_math_h_l739_c3_8d8d_return_output : unsigned(7 downto 0);

-- layer1_node2_MUX[bit_math_h_l750_c3_7ed6]
signal layer1_node2_MUX_bit_math_h_l750_c3_7ed6_cond : unsigned(0 downto 0);
signal layer1_node2_MUX_bit_math_h_l750_c3_7ed6_iftrue : unsigned(7 downto 0);
signal layer1_node2_MUX_bit_math_h_l750_c3_7ed6_iffalse : unsigned(7 downto 0);
signal layer1_node2_MUX_bit_math_h_l750_c3_7ed6_return_output : unsigned(7 downto 0);

-- layer1_node3_MUX[bit_math_h_l761_c3_68af]
signal layer1_node3_MUX_bit_math_h_l761_c3_68af_cond : unsigned(0 downto 0);
signal layer1_node3_MUX_bit_math_h_l761_c3_68af_iftrue : unsigned(7 downto 0);
signal layer1_node3_MUX_bit_math_h_l761_c3_68af_iffalse : unsigned(7 downto 0);
signal layer1_node3_MUX_bit_math_h_l761_c3_68af_return_output : unsigned(7 downto 0);

-- layer1_node4_MUX[bit_math_h_l772_c3_e8c5]
signal layer1_node4_MUX_bit_math_h_l772_c3_e8c5_cond : unsigned(0 downto 0);
signal layer1_node4_MUX_bit_math_h_l772_c3_e8c5_iftrue : unsigned(7 downto 0);
signal layer1_node4_MUX_bit_math_h_l772_c3_e8c5_iffalse : unsigned(7 downto 0);
signal layer1_node4_MUX_bit_math_h_l772_c3_e8c5_return_output : unsigned(7 downto 0);

-- layer1_node5_MUX[bit_math_h_l783_c3_7ab9]
signal layer1_node5_MUX_bit_math_h_l783_c3_7ab9_cond : unsigned(0 downto 0);
signal layer1_node5_MUX_bit_math_h_l783_c3_7ab9_iftrue : unsigned(7 downto 0);
signal layer1_node5_MUX_bit_math_h_l783_c3_7ab9_iffalse : unsigned(7 downto 0);
signal layer1_node5_MUX_bit_math_h_l783_c3_7ab9_return_output : unsigned(7 downto 0);

-- layer1_node6_MUX[bit_math_h_l794_c3_1dbe]
signal layer1_node6_MUX_bit_math_h_l794_c3_1dbe_cond : unsigned(0 downto 0);
signal layer1_node6_MUX_bit_math_h_l794_c3_1dbe_iftrue : unsigned(7 downto 0);
signal layer1_node6_MUX_bit_math_h_l794_c3_1dbe_iffalse : unsigned(7 downto 0);
signal layer1_node6_MUX_bit_math_h_l794_c3_1dbe_return_output : unsigned(7 downto 0);

-- layer1_node7_MUX[bit_math_h_l805_c3_6dfe]
signal layer1_node7_MUX_bit_math_h_l805_c3_6dfe_cond : unsigned(0 downto 0);
signal layer1_node7_MUX_bit_math_h_l805_c3_6dfe_iftrue : unsigned(7 downto 0);
signal layer1_node7_MUX_bit_math_h_l805_c3_6dfe_iffalse : unsigned(7 downto 0);
signal layer1_node7_MUX_bit_math_h_l805_c3_6dfe_return_output : unsigned(7 downto 0);

-- layer1_node8_MUX[bit_math_h_l816_c3_5d19]
signal layer1_node8_MUX_bit_math_h_l816_c3_5d19_cond : unsigned(0 downto 0);
signal layer1_node8_MUX_bit_math_h_l816_c3_5d19_iftrue : unsigned(7 downto 0);
signal layer1_node8_MUX_bit_math_h_l816_c3_5d19_iffalse : unsigned(7 downto 0);
signal layer1_node8_MUX_bit_math_h_l816_c3_5d19_return_output : unsigned(7 downto 0);

-- layer1_node9_MUX[bit_math_h_l827_c3_fe3d]
signal layer1_node9_MUX_bit_math_h_l827_c3_fe3d_cond : unsigned(0 downto 0);
signal layer1_node9_MUX_bit_math_h_l827_c3_fe3d_iftrue : unsigned(7 downto 0);
signal layer1_node9_MUX_bit_math_h_l827_c3_fe3d_iffalse : unsigned(7 downto 0);
signal layer1_node9_MUX_bit_math_h_l827_c3_fe3d_return_output : unsigned(7 downto 0);

-- layer1_node10_MUX[bit_math_h_l838_c3_cc59]
signal layer1_node10_MUX_bit_math_h_l838_c3_cc59_cond : unsigned(0 downto 0);
signal layer1_node10_MUX_bit_math_h_l838_c3_cc59_iftrue : unsigned(7 downto 0);
signal layer1_node10_MUX_bit_math_h_l838_c3_cc59_iffalse : unsigned(7 downto 0);
signal layer1_node10_MUX_bit_math_h_l838_c3_cc59_return_output : unsigned(7 downto 0);

-- layer1_node11_MUX[bit_math_h_l849_c3_6ba8]
signal layer1_node11_MUX_bit_math_h_l849_c3_6ba8_cond : unsigned(0 downto 0);
signal layer1_node11_MUX_bit_math_h_l849_c3_6ba8_iftrue : unsigned(7 downto 0);
signal layer1_node11_MUX_bit_math_h_l849_c3_6ba8_iffalse : unsigned(7 downto 0);
signal layer1_node11_MUX_bit_math_h_l849_c3_6ba8_return_output : unsigned(7 downto 0);

-- layer1_node12_MUX[bit_math_h_l860_c3_e057]
signal layer1_node12_MUX_bit_math_h_l860_c3_e057_cond : unsigned(0 downto 0);
signal layer1_node12_MUX_bit_math_h_l860_c3_e057_iftrue : unsigned(7 downto 0);
signal layer1_node12_MUX_bit_math_h_l860_c3_e057_iffalse : unsigned(7 downto 0);
signal layer1_node12_MUX_bit_math_h_l860_c3_e057_return_output : unsigned(7 downto 0);

-- layer1_node13_MUX[bit_math_h_l871_c3_aad3]
signal layer1_node13_MUX_bit_math_h_l871_c3_aad3_cond : unsigned(0 downto 0);
signal layer1_node13_MUX_bit_math_h_l871_c3_aad3_iftrue : unsigned(7 downto 0);
signal layer1_node13_MUX_bit_math_h_l871_c3_aad3_iffalse : unsigned(7 downto 0);
signal layer1_node13_MUX_bit_math_h_l871_c3_aad3_return_output : unsigned(7 downto 0);

-- layer1_node14_MUX[bit_math_h_l882_c3_0d3c]
signal layer1_node14_MUX_bit_math_h_l882_c3_0d3c_cond : unsigned(0 downto 0);
signal layer1_node14_MUX_bit_math_h_l882_c3_0d3c_iftrue : unsigned(7 downto 0);
signal layer1_node14_MUX_bit_math_h_l882_c3_0d3c_iffalse : unsigned(7 downto 0);
signal layer1_node14_MUX_bit_math_h_l882_c3_0d3c_return_output : unsigned(7 downto 0);

-- layer1_node15_MUX[bit_math_h_l893_c3_6301]
signal layer1_node15_MUX_bit_math_h_l893_c3_6301_cond : unsigned(0 downto 0);
signal layer1_node15_MUX_bit_math_h_l893_c3_6301_iftrue : unsigned(7 downto 0);
signal layer1_node15_MUX_bit_math_h_l893_c3_6301_iffalse : unsigned(7 downto 0);
signal layer1_node15_MUX_bit_math_h_l893_c3_6301_return_output : unsigned(7 downto 0);

-- layer1_node16_MUX[bit_math_h_l904_c3_60f0]
signal layer1_node16_MUX_bit_math_h_l904_c3_60f0_cond : unsigned(0 downto 0);
signal layer1_node16_MUX_bit_math_h_l904_c3_60f0_iftrue : unsigned(7 downto 0);
signal layer1_node16_MUX_bit_math_h_l904_c3_60f0_iffalse : unsigned(7 downto 0);
signal layer1_node16_MUX_bit_math_h_l904_c3_60f0_return_output : unsigned(7 downto 0);

-- layer1_node17_MUX[bit_math_h_l915_c3_d47f]
signal layer1_node17_MUX_bit_math_h_l915_c3_d47f_cond : unsigned(0 downto 0);
signal layer1_node17_MUX_bit_math_h_l915_c3_d47f_iftrue : unsigned(7 downto 0);
signal layer1_node17_MUX_bit_math_h_l915_c3_d47f_iffalse : unsigned(7 downto 0);
signal layer1_node17_MUX_bit_math_h_l915_c3_d47f_return_output : unsigned(7 downto 0);

-- layer1_node18_MUX[bit_math_h_l926_c3_678f]
signal layer1_node18_MUX_bit_math_h_l926_c3_678f_cond : unsigned(0 downto 0);
signal layer1_node18_MUX_bit_math_h_l926_c3_678f_iftrue : unsigned(7 downto 0);
signal layer1_node18_MUX_bit_math_h_l926_c3_678f_iffalse : unsigned(7 downto 0);
signal layer1_node18_MUX_bit_math_h_l926_c3_678f_return_output : unsigned(7 downto 0);

-- layer1_node19_MUX[bit_math_h_l937_c3_eb8f]
signal layer1_node19_MUX_bit_math_h_l937_c3_eb8f_cond : unsigned(0 downto 0);
signal layer1_node19_MUX_bit_math_h_l937_c3_eb8f_iftrue : unsigned(7 downto 0);
signal layer1_node19_MUX_bit_math_h_l937_c3_eb8f_iffalse : unsigned(7 downto 0);
signal layer1_node19_MUX_bit_math_h_l937_c3_eb8f_return_output : unsigned(7 downto 0);

-- layer1_node20_MUX[bit_math_h_l948_c3_588a]
signal layer1_node20_MUX_bit_math_h_l948_c3_588a_cond : unsigned(0 downto 0);
signal layer1_node20_MUX_bit_math_h_l948_c3_588a_iftrue : unsigned(7 downto 0);
signal layer1_node20_MUX_bit_math_h_l948_c3_588a_iffalse : unsigned(7 downto 0);
signal layer1_node20_MUX_bit_math_h_l948_c3_588a_return_output : unsigned(7 downto 0);

-- layer1_node21_MUX[bit_math_h_l959_c3_1823]
signal layer1_node21_MUX_bit_math_h_l959_c3_1823_cond : unsigned(0 downto 0);
signal layer1_node21_MUX_bit_math_h_l959_c3_1823_iftrue : unsigned(7 downto 0);
signal layer1_node21_MUX_bit_math_h_l959_c3_1823_iffalse : unsigned(7 downto 0);
signal layer1_node21_MUX_bit_math_h_l959_c3_1823_return_output : unsigned(7 downto 0);

-- layer1_node22_MUX[bit_math_h_l970_c3_6904]
signal layer1_node22_MUX_bit_math_h_l970_c3_6904_cond : unsigned(0 downto 0);
signal layer1_node22_MUX_bit_math_h_l970_c3_6904_iftrue : unsigned(7 downto 0);
signal layer1_node22_MUX_bit_math_h_l970_c3_6904_iffalse : unsigned(7 downto 0);
signal layer1_node22_MUX_bit_math_h_l970_c3_6904_return_output : unsigned(7 downto 0);

-- layer1_node23_MUX[bit_math_h_l981_c3_f890]
signal layer1_node23_MUX_bit_math_h_l981_c3_f890_cond : unsigned(0 downto 0);
signal layer1_node23_MUX_bit_math_h_l981_c3_f890_iftrue : unsigned(7 downto 0);
signal layer1_node23_MUX_bit_math_h_l981_c3_f890_iffalse : unsigned(7 downto 0);
signal layer1_node23_MUX_bit_math_h_l981_c3_f890_return_output : unsigned(7 downto 0);

-- layer1_node24_MUX[bit_math_h_l992_c3_4e65]
signal layer1_node24_MUX_bit_math_h_l992_c3_4e65_cond : unsigned(0 downto 0);
signal layer1_node24_MUX_bit_math_h_l992_c3_4e65_iftrue : unsigned(7 downto 0);
signal layer1_node24_MUX_bit_math_h_l992_c3_4e65_iffalse : unsigned(7 downto 0);
signal layer1_node24_MUX_bit_math_h_l992_c3_4e65_return_output : unsigned(7 downto 0);

-- layer1_node25_MUX[bit_math_h_l1003_c3_f943]
signal layer1_node25_MUX_bit_math_h_l1003_c3_f943_cond : unsigned(0 downto 0);
signal layer1_node25_MUX_bit_math_h_l1003_c3_f943_iftrue : unsigned(7 downto 0);
signal layer1_node25_MUX_bit_math_h_l1003_c3_f943_iffalse : unsigned(7 downto 0);
signal layer1_node25_MUX_bit_math_h_l1003_c3_f943_return_output : unsigned(7 downto 0);

-- layer1_node26_MUX[bit_math_h_l1014_c3_aa20]
signal layer1_node26_MUX_bit_math_h_l1014_c3_aa20_cond : unsigned(0 downto 0);
signal layer1_node26_MUX_bit_math_h_l1014_c3_aa20_iftrue : unsigned(7 downto 0);
signal layer1_node26_MUX_bit_math_h_l1014_c3_aa20_iffalse : unsigned(7 downto 0);
signal layer1_node26_MUX_bit_math_h_l1014_c3_aa20_return_output : unsigned(7 downto 0);

-- layer1_node27_MUX[bit_math_h_l1025_c3_a3a3]
signal layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_cond : unsigned(0 downto 0);
signal layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_iftrue : unsigned(7 downto 0);
signal layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_iffalse : unsigned(7 downto 0);
signal layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_return_output : unsigned(7 downto 0);

-- layer1_node28_MUX[bit_math_h_l1036_c3_85a0]
signal layer1_node28_MUX_bit_math_h_l1036_c3_85a0_cond : unsigned(0 downto 0);
signal layer1_node28_MUX_bit_math_h_l1036_c3_85a0_iftrue : unsigned(7 downto 0);
signal layer1_node28_MUX_bit_math_h_l1036_c3_85a0_iffalse : unsigned(7 downto 0);
signal layer1_node28_MUX_bit_math_h_l1036_c3_85a0_return_output : unsigned(7 downto 0);

-- layer1_node29_MUX[bit_math_h_l1047_c3_953f]
signal layer1_node29_MUX_bit_math_h_l1047_c3_953f_cond : unsigned(0 downto 0);
signal layer1_node29_MUX_bit_math_h_l1047_c3_953f_iftrue : unsigned(7 downto 0);
signal layer1_node29_MUX_bit_math_h_l1047_c3_953f_iffalse : unsigned(7 downto 0);
signal layer1_node29_MUX_bit_math_h_l1047_c3_953f_return_output : unsigned(7 downto 0);

-- layer1_node30_MUX[bit_math_h_l1058_c3_c3ba]
signal layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_cond : unsigned(0 downto 0);
signal layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_iftrue : unsigned(7 downto 0);
signal layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_iffalse : unsigned(7 downto 0);
signal layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_return_output : unsigned(7 downto 0);

-- layer1_node31_MUX[bit_math_h_l1069_c3_82fc]
signal layer1_node31_MUX_bit_math_h_l1069_c3_82fc_cond : unsigned(0 downto 0);
signal layer1_node31_MUX_bit_math_h_l1069_c3_82fc_iftrue : unsigned(7 downto 0);
signal layer1_node31_MUX_bit_math_h_l1069_c3_82fc_iffalse : unsigned(7 downto 0);
signal layer1_node31_MUX_bit_math_h_l1069_c3_82fc_return_output : unsigned(7 downto 0);

-- layer2_node0_MUX[bit_math_h_l1086_c3_4e60]
signal layer2_node0_MUX_bit_math_h_l1086_c3_4e60_cond : unsigned(0 downto 0);
signal layer2_node0_MUX_bit_math_h_l1086_c3_4e60_iftrue : unsigned(7 downto 0);
signal layer2_node0_MUX_bit_math_h_l1086_c3_4e60_iffalse : unsigned(7 downto 0);
signal layer2_node0_MUX_bit_math_h_l1086_c3_4e60_return_output : unsigned(7 downto 0);

-- layer2_node1_MUX[bit_math_h_l1097_c3_12bb]
signal layer2_node1_MUX_bit_math_h_l1097_c3_12bb_cond : unsigned(0 downto 0);
signal layer2_node1_MUX_bit_math_h_l1097_c3_12bb_iftrue : unsigned(7 downto 0);
signal layer2_node1_MUX_bit_math_h_l1097_c3_12bb_iffalse : unsigned(7 downto 0);
signal layer2_node1_MUX_bit_math_h_l1097_c3_12bb_return_output : unsigned(7 downto 0);

-- layer2_node2_MUX[bit_math_h_l1108_c3_fcbb]
signal layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_cond : unsigned(0 downto 0);
signal layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_iftrue : unsigned(7 downto 0);
signal layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_iffalse : unsigned(7 downto 0);
signal layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_return_output : unsigned(7 downto 0);

-- layer2_node3_MUX[bit_math_h_l1119_c3_8c7b]
signal layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_cond : unsigned(0 downto 0);
signal layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_iftrue : unsigned(7 downto 0);
signal layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_iffalse : unsigned(7 downto 0);
signal layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_return_output : unsigned(7 downto 0);

-- layer2_node4_MUX[bit_math_h_l1130_c3_3de0]
signal layer2_node4_MUX_bit_math_h_l1130_c3_3de0_cond : unsigned(0 downto 0);
signal layer2_node4_MUX_bit_math_h_l1130_c3_3de0_iftrue : unsigned(7 downto 0);
signal layer2_node4_MUX_bit_math_h_l1130_c3_3de0_iffalse : unsigned(7 downto 0);
signal layer2_node4_MUX_bit_math_h_l1130_c3_3de0_return_output : unsigned(7 downto 0);

-- layer2_node5_MUX[bit_math_h_l1141_c3_a5f6]
signal layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_cond : unsigned(0 downto 0);
signal layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_iftrue : unsigned(7 downto 0);
signal layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_iffalse : unsigned(7 downto 0);
signal layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_return_output : unsigned(7 downto 0);

-- layer2_node6_MUX[bit_math_h_l1152_c3_3828]
signal layer2_node6_MUX_bit_math_h_l1152_c3_3828_cond : unsigned(0 downto 0);
signal layer2_node6_MUX_bit_math_h_l1152_c3_3828_iftrue : unsigned(7 downto 0);
signal layer2_node6_MUX_bit_math_h_l1152_c3_3828_iffalse : unsigned(7 downto 0);
signal layer2_node6_MUX_bit_math_h_l1152_c3_3828_return_output : unsigned(7 downto 0);

-- layer2_node7_MUX[bit_math_h_l1163_c3_f226]
signal layer2_node7_MUX_bit_math_h_l1163_c3_f226_cond : unsigned(0 downto 0);
signal layer2_node7_MUX_bit_math_h_l1163_c3_f226_iftrue : unsigned(7 downto 0);
signal layer2_node7_MUX_bit_math_h_l1163_c3_f226_iffalse : unsigned(7 downto 0);
signal layer2_node7_MUX_bit_math_h_l1163_c3_f226_return_output : unsigned(7 downto 0);

-- layer2_node8_MUX[bit_math_h_l1174_c3_49b7]
signal layer2_node8_MUX_bit_math_h_l1174_c3_49b7_cond : unsigned(0 downto 0);
signal layer2_node8_MUX_bit_math_h_l1174_c3_49b7_iftrue : unsigned(7 downto 0);
signal layer2_node8_MUX_bit_math_h_l1174_c3_49b7_iffalse : unsigned(7 downto 0);
signal layer2_node8_MUX_bit_math_h_l1174_c3_49b7_return_output : unsigned(7 downto 0);

-- layer2_node9_MUX[bit_math_h_l1185_c3_934f]
signal layer2_node9_MUX_bit_math_h_l1185_c3_934f_cond : unsigned(0 downto 0);
signal layer2_node9_MUX_bit_math_h_l1185_c3_934f_iftrue : unsigned(7 downto 0);
signal layer2_node9_MUX_bit_math_h_l1185_c3_934f_iffalse : unsigned(7 downto 0);
signal layer2_node9_MUX_bit_math_h_l1185_c3_934f_return_output : unsigned(7 downto 0);

-- layer2_node10_MUX[bit_math_h_l1196_c3_3f7c]
signal layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_cond : unsigned(0 downto 0);
signal layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_iftrue : unsigned(7 downto 0);
signal layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_iffalse : unsigned(7 downto 0);
signal layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_return_output : unsigned(7 downto 0);

-- layer2_node11_MUX[bit_math_h_l1207_c3_d0a7]
signal layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_cond : unsigned(0 downto 0);
signal layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_iftrue : unsigned(7 downto 0);
signal layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_iffalse : unsigned(7 downto 0);
signal layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_return_output : unsigned(7 downto 0);

-- layer2_node12_MUX[bit_math_h_l1218_c3_0726]
signal layer2_node12_MUX_bit_math_h_l1218_c3_0726_cond : unsigned(0 downto 0);
signal layer2_node12_MUX_bit_math_h_l1218_c3_0726_iftrue : unsigned(7 downto 0);
signal layer2_node12_MUX_bit_math_h_l1218_c3_0726_iffalse : unsigned(7 downto 0);
signal layer2_node12_MUX_bit_math_h_l1218_c3_0726_return_output : unsigned(7 downto 0);

-- layer2_node13_MUX[bit_math_h_l1229_c3_754d]
signal layer2_node13_MUX_bit_math_h_l1229_c3_754d_cond : unsigned(0 downto 0);
signal layer2_node13_MUX_bit_math_h_l1229_c3_754d_iftrue : unsigned(7 downto 0);
signal layer2_node13_MUX_bit_math_h_l1229_c3_754d_iffalse : unsigned(7 downto 0);
signal layer2_node13_MUX_bit_math_h_l1229_c3_754d_return_output : unsigned(7 downto 0);

-- layer2_node14_MUX[bit_math_h_l1240_c3_2b9a]
signal layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_cond : unsigned(0 downto 0);
signal layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_iftrue : unsigned(7 downto 0);
signal layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_iffalse : unsigned(7 downto 0);
signal layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_return_output : unsigned(7 downto 0);

-- layer2_node15_MUX[bit_math_h_l1251_c3_57b2]
signal layer2_node15_MUX_bit_math_h_l1251_c3_57b2_cond : unsigned(0 downto 0);
signal layer2_node15_MUX_bit_math_h_l1251_c3_57b2_iftrue : unsigned(7 downto 0);
signal layer2_node15_MUX_bit_math_h_l1251_c3_57b2_iffalse : unsigned(7 downto 0);
signal layer2_node15_MUX_bit_math_h_l1251_c3_57b2_return_output : unsigned(7 downto 0);

-- layer3_node0_MUX[bit_math_h_l1268_c3_e5cc]
signal layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_cond : unsigned(0 downto 0);
signal layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_iftrue : unsigned(7 downto 0);
signal layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_iffalse : unsigned(7 downto 0);
signal layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_return_output : unsigned(7 downto 0);

-- layer3_node1_MUX[bit_math_h_l1279_c3_73ae]
signal layer3_node1_MUX_bit_math_h_l1279_c3_73ae_cond : unsigned(0 downto 0);
signal layer3_node1_MUX_bit_math_h_l1279_c3_73ae_iftrue : unsigned(7 downto 0);
signal layer3_node1_MUX_bit_math_h_l1279_c3_73ae_iffalse : unsigned(7 downto 0);
signal layer3_node1_MUX_bit_math_h_l1279_c3_73ae_return_output : unsigned(7 downto 0);

-- layer3_node2_MUX[bit_math_h_l1290_c3_d8d2]
signal layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_cond : unsigned(0 downto 0);
signal layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_iftrue : unsigned(7 downto 0);
signal layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_iffalse : unsigned(7 downto 0);
signal layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_return_output : unsigned(7 downto 0);

-- layer3_node3_MUX[bit_math_h_l1301_c3_827d]
signal layer3_node3_MUX_bit_math_h_l1301_c3_827d_cond : unsigned(0 downto 0);
signal layer3_node3_MUX_bit_math_h_l1301_c3_827d_iftrue : unsigned(7 downto 0);
signal layer3_node3_MUX_bit_math_h_l1301_c3_827d_iffalse : unsigned(7 downto 0);
signal layer3_node3_MUX_bit_math_h_l1301_c3_827d_return_output : unsigned(7 downto 0);

-- layer3_node4_MUX[bit_math_h_l1312_c3_ca04]
signal layer3_node4_MUX_bit_math_h_l1312_c3_ca04_cond : unsigned(0 downto 0);
signal layer3_node4_MUX_bit_math_h_l1312_c3_ca04_iftrue : unsigned(7 downto 0);
signal layer3_node4_MUX_bit_math_h_l1312_c3_ca04_iffalse : unsigned(7 downto 0);
signal layer3_node4_MUX_bit_math_h_l1312_c3_ca04_return_output : unsigned(7 downto 0);

-- layer3_node5_MUX[bit_math_h_l1323_c3_56dd]
signal layer3_node5_MUX_bit_math_h_l1323_c3_56dd_cond : unsigned(0 downto 0);
signal layer3_node5_MUX_bit_math_h_l1323_c3_56dd_iftrue : unsigned(7 downto 0);
signal layer3_node5_MUX_bit_math_h_l1323_c3_56dd_iffalse : unsigned(7 downto 0);
signal layer3_node5_MUX_bit_math_h_l1323_c3_56dd_return_output : unsigned(7 downto 0);

-- layer3_node6_MUX[bit_math_h_l1334_c3_07bd]
signal layer3_node6_MUX_bit_math_h_l1334_c3_07bd_cond : unsigned(0 downto 0);
signal layer3_node6_MUX_bit_math_h_l1334_c3_07bd_iftrue : unsigned(7 downto 0);
signal layer3_node6_MUX_bit_math_h_l1334_c3_07bd_iffalse : unsigned(7 downto 0);
signal layer3_node6_MUX_bit_math_h_l1334_c3_07bd_return_output : unsigned(7 downto 0);

-- layer3_node7_MUX[bit_math_h_l1345_c3_5a50]
signal layer3_node7_MUX_bit_math_h_l1345_c3_5a50_cond : unsigned(0 downto 0);
signal layer3_node7_MUX_bit_math_h_l1345_c3_5a50_iftrue : unsigned(7 downto 0);
signal layer3_node7_MUX_bit_math_h_l1345_c3_5a50_iffalse : unsigned(7 downto 0);
signal layer3_node7_MUX_bit_math_h_l1345_c3_5a50_return_output : unsigned(7 downto 0);

-- layer4_node0_MUX[bit_math_h_l1362_c3_f5a3]
signal layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_cond : unsigned(0 downto 0);
signal layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_iftrue : unsigned(7 downto 0);
signal layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_iffalse : unsigned(7 downto 0);
signal layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_return_output : unsigned(7 downto 0);

-- layer4_node1_MUX[bit_math_h_l1373_c3_402b]
signal layer4_node1_MUX_bit_math_h_l1373_c3_402b_cond : unsigned(0 downto 0);
signal layer4_node1_MUX_bit_math_h_l1373_c3_402b_iftrue : unsigned(7 downto 0);
signal layer4_node1_MUX_bit_math_h_l1373_c3_402b_iffalse : unsigned(7 downto 0);
signal layer4_node1_MUX_bit_math_h_l1373_c3_402b_return_output : unsigned(7 downto 0);

-- layer4_node2_MUX[bit_math_h_l1384_c3_5f80]
signal layer4_node2_MUX_bit_math_h_l1384_c3_5f80_cond : unsigned(0 downto 0);
signal layer4_node2_MUX_bit_math_h_l1384_c3_5f80_iftrue : unsigned(7 downto 0);
signal layer4_node2_MUX_bit_math_h_l1384_c3_5f80_iffalse : unsigned(7 downto 0);
signal layer4_node2_MUX_bit_math_h_l1384_c3_5f80_return_output : unsigned(7 downto 0);

-- layer4_node3_MUX[bit_math_h_l1395_c3_4d9c]
signal layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_cond : unsigned(0 downto 0);
signal layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_iftrue : unsigned(7 downto 0);
signal layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_iffalse : unsigned(7 downto 0);
signal layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_return_output : unsigned(7 downto 0);

-- layer5_node0_MUX[bit_math_h_l1412_c3_19e3]
signal layer5_node0_MUX_bit_math_h_l1412_c3_19e3_cond : unsigned(0 downto 0);
signal layer5_node0_MUX_bit_math_h_l1412_c3_19e3_iftrue : unsigned(7 downto 0);
signal layer5_node0_MUX_bit_math_h_l1412_c3_19e3_iffalse : unsigned(7 downto 0);
signal layer5_node0_MUX_bit_math_h_l1412_c3_19e3_return_output : unsigned(7 downto 0);

-- layer5_node1_MUX[bit_math_h_l1423_c3_11f1]
signal layer5_node1_MUX_bit_math_h_l1423_c3_11f1_cond : unsigned(0 downto 0);
signal layer5_node1_MUX_bit_math_h_l1423_c3_11f1_iftrue : unsigned(7 downto 0);
signal layer5_node1_MUX_bit_math_h_l1423_c3_11f1_iffalse : unsigned(7 downto 0);
signal layer5_node1_MUX_bit_math_h_l1423_c3_11f1_return_output : unsigned(7 downto 0);

-- layer6_node0_MUX[bit_math_h_l1440_c3_f906]
signal layer6_node0_MUX_bit_math_h_l1440_c3_f906_cond : unsigned(0 downto 0);
signal layer6_node0_MUX_bit_math_h_l1440_c3_f906_iftrue : unsigned(7 downto 0);
signal layer6_node0_MUX_bit_math_h_l1440_c3_f906_iffalse : unsigned(7 downto 0);
signal layer6_node0_MUX_bit_math_h_l1440_c3_f906_return_output : unsigned(7 downto 0);

function uint7_0_0( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(0- i);
      end loop;
return return_output;
end function;

function uint7_1_1( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(1- i);
      end loop;
return return_output;
end function;

function uint7_2_2( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(2- i);
      end loop;
return return_output;
end function;

function uint7_3_3( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(3- i);
      end loop;
return return_output;
end function;

function uint7_4_4( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(4- i);
      end loop;
return return_output;
end function;

function uint7_5_5( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(5- i);
      end loop;
return return_output;
end function;

function uint7_6_6( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(6- i);
      end loop;
return return_output;
end function;


begin

-- SUBMODULE INSTANCES 
-- layer0_node0_MUX_bit_math_h_l18_c3_5c06
layer0_node0_MUX_bit_math_h_l18_c3_5c06 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node0_MUX_bit_math_h_l18_c3_5c06_cond,
layer0_node0_MUX_bit_math_h_l18_c3_5c06_iftrue,
layer0_node0_MUX_bit_math_h_l18_c3_5c06_iffalse,
layer0_node0_MUX_bit_math_h_l18_c3_5c06_return_output);

-- layer0_node1_MUX_bit_math_h_l29_c3_fa46
layer0_node1_MUX_bit_math_h_l29_c3_fa46 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node1_MUX_bit_math_h_l29_c3_fa46_cond,
layer0_node1_MUX_bit_math_h_l29_c3_fa46_iftrue,
layer0_node1_MUX_bit_math_h_l29_c3_fa46_iffalse,
layer0_node1_MUX_bit_math_h_l29_c3_fa46_return_output);

-- layer0_node2_MUX_bit_math_h_l40_c3_f68a
layer0_node2_MUX_bit_math_h_l40_c3_f68a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node2_MUX_bit_math_h_l40_c3_f68a_cond,
layer0_node2_MUX_bit_math_h_l40_c3_f68a_iftrue,
layer0_node2_MUX_bit_math_h_l40_c3_f68a_iffalse,
layer0_node2_MUX_bit_math_h_l40_c3_f68a_return_output);

-- layer0_node3_MUX_bit_math_h_l51_c3_b336
layer0_node3_MUX_bit_math_h_l51_c3_b336 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node3_MUX_bit_math_h_l51_c3_b336_cond,
layer0_node3_MUX_bit_math_h_l51_c3_b336_iftrue,
layer0_node3_MUX_bit_math_h_l51_c3_b336_iffalse,
layer0_node3_MUX_bit_math_h_l51_c3_b336_return_output);

-- layer0_node4_MUX_bit_math_h_l62_c3_07e7
layer0_node4_MUX_bit_math_h_l62_c3_07e7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node4_MUX_bit_math_h_l62_c3_07e7_cond,
layer0_node4_MUX_bit_math_h_l62_c3_07e7_iftrue,
layer0_node4_MUX_bit_math_h_l62_c3_07e7_iffalse,
layer0_node4_MUX_bit_math_h_l62_c3_07e7_return_output);

-- layer0_node5_MUX_bit_math_h_l73_c3_282b
layer0_node5_MUX_bit_math_h_l73_c3_282b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node5_MUX_bit_math_h_l73_c3_282b_cond,
layer0_node5_MUX_bit_math_h_l73_c3_282b_iftrue,
layer0_node5_MUX_bit_math_h_l73_c3_282b_iffalse,
layer0_node5_MUX_bit_math_h_l73_c3_282b_return_output);

-- layer0_node6_MUX_bit_math_h_l84_c3_62f1
layer0_node6_MUX_bit_math_h_l84_c3_62f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node6_MUX_bit_math_h_l84_c3_62f1_cond,
layer0_node6_MUX_bit_math_h_l84_c3_62f1_iftrue,
layer0_node6_MUX_bit_math_h_l84_c3_62f1_iffalse,
layer0_node6_MUX_bit_math_h_l84_c3_62f1_return_output);

-- layer0_node7_MUX_bit_math_h_l95_c3_567b
layer0_node7_MUX_bit_math_h_l95_c3_567b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node7_MUX_bit_math_h_l95_c3_567b_cond,
layer0_node7_MUX_bit_math_h_l95_c3_567b_iftrue,
layer0_node7_MUX_bit_math_h_l95_c3_567b_iffalse,
layer0_node7_MUX_bit_math_h_l95_c3_567b_return_output);

-- layer0_node8_MUX_bit_math_h_l106_c3_47e5
layer0_node8_MUX_bit_math_h_l106_c3_47e5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node8_MUX_bit_math_h_l106_c3_47e5_cond,
layer0_node8_MUX_bit_math_h_l106_c3_47e5_iftrue,
layer0_node8_MUX_bit_math_h_l106_c3_47e5_iffalse,
layer0_node8_MUX_bit_math_h_l106_c3_47e5_return_output);

-- layer0_node9_MUX_bit_math_h_l117_c3_f097
layer0_node9_MUX_bit_math_h_l117_c3_f097 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node9_MUX_bit_math_h_l117_c3_f097_cond,
layer0_node9_MUX_bit_math_h_l117_c3_f097_iftrue,
layer0_node9_MUX_bit_math_h_l117_c3_f097_iffalse,
layer0_node9_MUX_bit_math_h_l117_c3_f097_return_output);

-- layer0_node10_MUX_bit_math_h_l128_c3_0e6c
layer0_node10_MUX_bit_math_h_l128_c3_0e6c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node10_MUX_bit_math_h_l128_c3_0e6c_cond,
layer0_node10_MUX_bit_math_h_l128_c3_0e6c_iftrue,
layer0_node10_MUX_bit_math_h_l128_c3_0e6c_iffalse,
layer0_node10_MUX_bit_math_h_l128_c3_0e6c_return_output);

-- layer0_node11_MUX_bit_math_h_l139_c3_3ab9
layer0_node11_MUX_bit_math_h_l139_c3_3ab9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node11_MUX_bit_math_h_l139_c3_3ab9_cond,
layer0_node11_MUX_bit_math_h_l139_c3_3ab9_iftrue,
layer0_node11_MUX_bit_math_h_l139_c3_3ab9_iffalse,
layer0_node11_MUX_bit_math_h_l139_c3_3ab9_return_output);

-- layer0_node12_MUX_bit_math_h_l150_c3_e611
layer0_node12_MUX_bit_math_h_l150_c3_e611 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node12_MUX_bit_math_h_l150_c3_e611_cond,
layer0_node12_MUX_bit_math_h_l150_c3_e611_iftrue,
layer0_node12_MUX_bit_math_h_l150_c3_e611_iffalse,
layer0_node12_MUX_bit_math_h_l150_c3_e611_return_output);

-- layer0_node13_MUX_bit_math_h_l161_c3_e037
layer0_node13_MUX_bit_math_h_l161_c3_e037 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node13_MUX_bit_math_h_l161_c3_e037_cond,
layer0_node13_MUX_bit_math_h_l161_c3_e037_iftrue,
layer0_node13_MUX_bit_math_h_l161_c3_e037_iffalse,
layer0_node13_MUX_bit_math_h_l161_c3_e037_return_output);

-- layer0_node14_MUX_bit_math_h_l172_c3_ad25
layer0_node14_MUX_bit_math_h_l172_c3_ad25 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node14_MUX_bit_math_h_l172_c3_ad25_cond,
layer0_node14_MUX_bit_math_h_l172_c3_ad25_iftrue,
layer0_node14_MUX_bit_math_h_l172_c3_ad25_iffalse,
layer0_node14_MUX_bit_math_h_l172_c3_ad25_return_output);

-- layer0_node15_MUX_bit_math_h_l183_c3_dacd
layer0_node15_MUX_bit_math_h_l183_c3_dacd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node15_MUX_bit_math_h_l183_c3_dacd_cond,
layer0_node15_MUX_bit_math_h_l183_c3_dacd_iftrue,
layer0_node15_MUX_bit_math_h_l183_c3_dacd_iffalse,
layer0_node15_MUX_bit_math_h_l183_c3_dacd_return_output);

-- layer0_node16_MUX_bit_math_h_l194_c3_5393
layer0_node16_MUX_bit_math_h_l194_c3_5393 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node16_MUX_bit_math_h_l194_c3_5393_cond,
layer0_node16_MUX_bit_math_h_l194_c3_5393_iftrue,
layer0_node16_MUX_bit_math_h_l194_c3_5393_iffalse,
layer0_node16_MUX_bit_math_h_l194_c3_5393_return_output);

-- layer0_node17_MUX_bit_math_h_l205_c3_4246
layer0_node17_MUX_bit_math_h_l205_c3_4246 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node17_MUX_bit_math_h_l205_c3_4246_cond,
layer0_node17_MUX_bit_math_h_l205_c3_4246_iftrue,
layer0_node17_MUX_bit_math_h_l205_c3_4246_iffalse,
layer0_node17_MUX_bit_math_h_l205_c3_4246_return_output);

-- layer0_node18_MUX_bit_math_h_l216_c3_2748
layer0_node18_MUX_bit_math_h_l216_c3_2748 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node18_MUX_bit_math_h_l216_c3_2748_cond,
layer0_node18_MUX_bit_math_h_l216_c3_2748_iftrue,
layer0_node18_MUX_bit_math_h_l216_c3_2748_iffalse,
layer0_node18_MUX_bit_math_h_l216_c3_2748_return_output);

-- layer0_node19_MUX_bit_math_h_l227_c3_1dae
layer0_node19_MUX_bit_math_h_l227_c3_1dae : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node19_MUX_bit_math_h_l227_c3_1dae_cond,
layer0_node19_MUX_bit_math_h_l227_c3_1dae_iftrue,
layer0_node19_MUX_bit_math_h_l227_c3_1dae_iffalse,
layer0_node19_MUX_bit_math_h_l227_c3_1dae_return_output);

-- layer0_node20_MUX_bit_math_h_l238_c3_e7c7
layer0_node20_MUX_bit_math_h_l238_c3_e7c7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node20_MUX_bit_math_h_l238_c3_e7c7_cond,
layer0_node20_MUX_bit_math_h_l238_c3_e7c7_iftrue,
layer0_node20_MUX_bit_math_h_l238_c3_e7c7_iffalse,
layer0_node20_MUX_bit_math_h_l238_c3_e7c7_return_output);

-- layer0_node21_MUX_bit_math_h_l249_c3_8f8c
layer0_node21_MUX_bit_math_h_l249_c3_8f8c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node21_MUX_bit_math_h_l249_c3_8f8c_cond,
layer0_node21_MUX_bit_math_h_l249_c3_8f8c_iftrue,
layer0_node21_MUX_bit_math_h_l249_c3_8f8c_iffalse,
layer0_node21_MUX_bit_math_h_l249_c3_8f8c_return_output);

-- layer0_node22_MUX_bit_math_h_l260_c3_321e
layer0_node22_MUX_bit_math_h_l260_c3_321e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node22_MUX_bit_math_h_l260_c3_321e_cond,
layer0_node22_MUX_bit_math_h_l260_c3_321e_iftrue,
layer0_node22_MUX_bit_math_h_l260_c3_321e_iffalse,
layer0_node22_MUX_bit_math_h_l260_c3_321e_return_output);

-- layer0_node23_MUX_bit_math_h_l271_c3_86c3
layer0_node23_MUX_bit_math_h_l271_c3_86c3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node23_MUX_bit_math_h_l271_c3_86c3_cond,
layer0_node23_MUX_bit_math_h_l271_c3_86c3_iftrue,
layer0_node23_MUX_bit_math_h_l271_c3_86c3_iffalse,
layer0_node23_MUX_bit_math_h_l271_c3_86c3_return_output);

-- layer0_node24_MUX_bit_math_h_l282_c3_2992
layer0_node24_MUX_bit_math_h_l282_c3_2992 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node24_MUX_bit_math_h_l282_c3_2992_cond,
layer0_node24_MUX_bit_math_h_l282_c3_2992_iftrue,
layer0_node24_MUX_bit_math_h_l282_c3_2992_iffalse,
layer0_node24_MUX_bit_math_h_l282_c3_2992_return_output);

-- layer0_node25_MUX_bit_math_h_l293_c3_ece2
layer0_node25_MUX_bit_math_h_l293_c3_ece2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node25_MUX_bit_math_h_l293_c3_ece2_cond,
layer0_node25_MUX_bit_math_h_l293_c3_ece2_iftrue,
layer0_node25_MUX_bit_math_h_l293_c3_ece2_iffalse,
layer0_node25_MUX_bit_math_h_l293_c3_ece2_return_output);

-- layer0_node26_MUX_bit_math_h_l304_c3_7f9b
layer0_node26_MUX_bit_math_h_l304_c3_7f9b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node26_MUX_bit_math_h_l304_c3_7f9b_cond,
layer0_node26_MUX_bit_math_h_l304_c3_7f9b_iftrue,
layer0_node26_MUX_bit_math_h_l304_c3_7f9b_iffalse,
layer0_node26_MUX_bit_math_h_l304_c3_7f9b_return_output);

-- layer0_node27_MUX_bit_math_h_l315_c3_5c0f
layer0_node27_MUX_bit_math_h_l315_c3_5c0f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node27_MUX_bit_math_h_l315_c3_5c0f_cond,
layer0_node27_MUX_bit_math_h_l315_c3_5c0f_iftrue,
layer0_node27_MUX_bit_math_h_l315_c3_5c0f_iffalse,
layer0_node27_MUX_bit_math_h_l315_c3_5c0f_return_output);

-- layer0_node28_MUX_bit_math_h_l326_c3_12a3
layer0_node28_MUX_bit_math_h_l326_c3_12a3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node28_MUX_bit_math_h_l326_c3_12a3_cond,
layer0_node28_MUX_bit_math_h_l326_c3_12a3_iftrue,
layer0_node28_MUX_bit_math_h_l326_c3_12a3_iffalse,
layer0_node28_MUX_bit_math_h_l326_c3_12a3_return_output);

-- layer0_node29_MUX_bit_math_h_l337_c3_cbb8
layer0_node29_MUX_bit_math_h_l337_c3_cbb8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node29_MUX_bit_math_h_l337_c3_cbb8_cond,
layer0_node29_MUX_bit_math_h_l337_c3_cbb8_iftrue,
layer0_node29_MUX_bit_math_h_l337_c3_cbb8_iffalse,
layer0_node29_MUX_bit_math_h_l337_c3_cbb8_return_output);

-- layer0_node30_MUX_bit_math_h_l348_c3_8c5c
layer0_node30_MUX_bit_math_h_l348_c3_8c5c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node30_MUX_bit_math_h_l348_c3_8c5c_cond,
layer0_node30_MUX_bit_math_h_l348_c3_8c5c_iftrue,
layer0_node30_MUX_bit_math_h_l348_c3_8c5c_iffalse,
layer0_node30_MUX_bit_math_h_l348_c3_8c5c_return_output);

-- layer0_node31_MUX_bit_math_h_l359_c3_d6b9
layer0_node31_MUX_bit_math_h_l359_c3_d6b9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node31_MUX_bit_math_h_l359_c3_d6b9_cond,
layer0_node31_MUX_bit_math_h_l359_c3_d6b9_iftrue,
layer0_node31_MUX_bit_math_h_l359_c3_d6b9_iffalse,
layer0_node31_MUX_bit_math_h_l359_c3_d6b9_return_output);

-- layer0_node32_MUX_bit_math_h_l370_c3_3d24
layer0_node32_MUX_bit_math_h_l370_c3_3d24 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node32_MUX_bit_math_h_l370_c3_3d24_cond,
layer0_node32_MUX_bit_math_h_l370_c3_3d24_iftrue,
layer0_node32_MUX_bit_math_h_l370_c3_3d24_iffalse,
layer0_node32_MUX_bit_math_h_l370_c3_3d24_return_output);

-- layer0_node33_MUX_bit_math_h_l381_c3_bdd0
layer0_node33_MUX_bit_math_h_l381_c3_bdd0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node33_MUX_bit_math_h_l381_c3_bdd0_cond,
layer0_node33_MUX_bit_math_h_l381_c3_bdd0_iftrue,
layer0_node33_MUX_bit_math_h_l381_c3_bdd0_iffalse,
layer0_node33_MUX_bit_math_h_l381_c3_bdd0_return_output);

-- layer0_node34_MUX_bit_math_h_l392_c3_f617
layer0_node34_MUX_bit_math_h_l392_c3_f617 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node34_MUX_bit_math_h_l392_c3_f617_cond,
layer0_node34_MUX_bit_math_h_l392_c3_f617_iftrue,
layer0_node34_MUX_bit_math_h_l392_c3_f617_iffalse,
layer0_node34_MUX_bit_math_h_l392_c3_f617_return_output);

-- layer0_node35_MUX_bit_math_h_l403_c3_683e
layer0_node35_MUX_bit_math_h_l403_c3_683e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node35_MUX_bit_math_h_l403_c3_683e_cond,
layer0_node35_MUX_bit_math_h_l403_c3_683e_iftrue,
layer0_node35_MUX_bit_math_h_l403_c3_683e_iffalse,
layer0_node35_MUX_bit_math_h_l403_c3_683e_return_output);

-- layer0_node36_MUX_bit_math_h_l414_c3_cd2c
layer0_node36_MUX_bit_math_h_l414_c3_cd2c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node36_MUX_bit_math_h_l414_c3_cd2c_cond,
layer0_node36_MUX_bit_math_h_l414_c3_cd2c_iftrue,
layer0_node36_MUX_bit_math_h_l414_c3_cd2c_iffalse,
layer0_node36_MUX_bit_math_h_l414_c3_cd2c_return_output);

-- layer0_node37_MUX_bit_math_h_l425_c3_2485
layer0_node37_MUX_bit_math_h_l425_c3_2485 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node37_MUX_bit_math_h_l425_c3_2485_cond,
layer0_node37_MUX_bit_math_h_l425_c3_2485_iftrue,
layer0_node37_MUX_bit_math_h_l425_c3_2485_iffalse,
layer0_node37_MUX_bit_math_h_l425_c3_2485_return_output);

-- layer0_node38_MUX_bit_math_h_l436_c3_c940
layer0_node38_MUX_bit_math_h_l436_c3_c940 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node38_MUX_bit_math_h_l436_c3_c940_cond,
layer0_node38_MUX_bit_math_h_l436_c3_c940_iftrue,
layer0_node38_MUX_bit_math_h_l436_c3_c940_iffalse,
layer0_node38_MUX_bit_math_h_l436_c3_c940_return_output);

-- layer0_node39_MUX_bit_math_h_l447_c3_b150
layer0_node39_MUX_bit_math_h_l447_c3_b150 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node39_MUX_bit_math_h_l447_c3_b150_cond,
layer0_node39_MUX_bit_math_h_l447_c3_b150_iftrue,
layer0_node39_MUX_bit_math_h_l447_c3_b150_iffalse,
layer0_node39_MUX_bit_math_h_l447_c3_b150_return_output);

-- layer0_node40_MUX_bit_math_h_l458_c3_c977
layer0_node40_MUX_bit_math_h_l458_c3_c977 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node40_MUX_bit_math_h_l458_c3_c977_cond,
layer0_node40_MUX_bit_math_h_l458_c3_c977_iftrue,
layer0_node40_MUX_bit_math_h_l458_c3_c977_iffalse,
layer0_node40_MUX_bit_math_h_l458_c3_c977_return_output);

-- layer0_node41_MUX_bit_math_h_l469_c3_b3bf
layer0_node41_MUX_bit_math_h_l469_c3_b3bf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node41_MUX_bit_math_h_l469_c3_b3bf_cond,
layer0_node41_MUX_bit_math_h_l469_c3_b3bf_iftrue,
layer0_node41_MUX_bit_math_h_l469_c3_b3bf_iffalse,
layer0_node41_MUX_bit_math_h_l469_c3_b3bf_return_output);

-- layer0_node42_MUX_bit_math_h_l480_c3_c677
layer0_node42_MUX_bit_math_h_l480_c3_c677 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node42_MUX_bit_math_h_l480_c3_c677_cond,
layer0_node42_MUX_bit_math_h_l480_c3_c677_iftrue,
layer0_node42_MUX_bit_math_h_l480_c3_c677_iffalse,
layer0_node42_MUX_bit_math_h_l480_c3_c677_return_output);

-- layer0_node43_MUX_bit_math_h_l491_c3_2838
layer0_node43_MUX_bit_math_h_l491_c3_2838 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node43_MUX_bit_math_h_l491_c3_2838_cond,
layer0_node43_MUX_bit_math_h_l491_c3_2838_iftrue,
layer0_node43_MUX_bit_math_h_l491_c3_2838_iffalse,
layer0_node43_MUX_bit_math_h_l491_c3_2838_return_output);

-- layer0_node44_MUX_bit_math_h_l502_c3_6b96
layer0_node44_MUX_bit_math_h_l502_c3_6b96 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node44_MUX_bit_math_h_l502_c3_6b96_cond,
layer0_node44_MUX_bit_math_h_l502_c3_6b96_iftrue,
layer0_node44_MUX_bit_math_h_l502_c3_6b96_iffalse,
layer0_node44_MUX_bit_math_h_l502_c3_6b96_return_output);

-- layer0_node45_MUX_bit_math_h_l513_c3_b86e
layer0_node45_MUX_bit_math_h_l513_c3_b86e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node45_MUX_bit_math_h_l513_c3_b86e_cond,
layer0_node45_MUX_bit_math_h_l513_c3_b86e_iftrue,
layer0_node45_MUX_bit_math_h_l513_c3_b86e_iffalse,
layer0_node45_MUX_bit_math_h_l513_c3_b86e_return_output);

-- layer0_node46_MUX_bit_math_h_l524_c3_4ef5
layer0_node46_MUX_bit_math_h_l524_c3_4ef5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node46_MUX_bit_math_h_l524_c3_4ef5_cond,
layer0_node46_MUX_bit_math_h_l524_c3_4ef5_iftrue,
layer0_node46_MUX_bit_math_h_l524_c3_4ef5_iffalse,
layer0_node46_MUX_bit_math_h_l524_c3_4ef5_return_output);

-- layer0_node47_MUX_bit_math_h_l535_c3_21f3
layer0_node47_MUX_bit_math_h_l535_c3_21f3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node47_MUX_bit_math_h_l535_c3_21f3_cond,
layer0_node47_MUX_bit_math_h_l535_c3_21f3_iftrue,
layer0_node47_MUX_bit_math_h_l535_c3_21f3_iffalse,
layer0_node47_MUX_bit_math_h_l535_c3_21f3_return_output);

-- layer0_node48_MUX_bit_math_h_l546_c3_5be4
layer0_node48_MUX_bit_math_h_l546_c3_5be4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node48_MUX_bit_math_h_l546_c3_5be4_cond,
layer0_node48_MUX_bit_math_h_l546_c3_5be4_iftrue,
layer0_node48_MUX_bit_math_h_l546_c3_5be4_iffalse,
layer0_node48_MUX_bit_math_h_l546_c3_5be4_return_output);

-- layer0_node49_MUX_bit_math_h_l557_c3_3410
layer0_node49_MUX_bit_math_h_l557_c3_3410 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node49_MUX_bit_math_h_l557_c3_3410_cond,
layer0_node49_MUX_bit_math_h_l557_c3_3410_iftrue,
layer0_node49_MUX_bit_math_h_l557_c3_3410_iffalse,
layer0_node49_MUX_bit_math_h_l557_c3_3410_return_output);

-- layer0_node50_MUX_bit_math_h_l568_c3_4522
layer0_node50_MUX_bit_math_h_l568_c3_4522 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node50_MUX_bit_math_h_l568_c3_4522_cond,
layer0_node50_MUX_bit_math_h_l568_c3_4522_iftrue,
layer0_node50_MUX_bit_math_h_l568_c3_4522_iffalse,
layer0_node50_MUX_bit_math_h_l568_c3_4522_return_output);

-- layer0_node51_MUX_bit_math_h_l579_c3_8398
layer0_node51_MUX_bit_math_h_l579_c3_8398 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node51_MUX_bit_math_h_l579_c3_8398_cond,
layer0_node51_MUX_bit_math_h_l579_c3_8398_iftrue,
layer0_node51_MUX_bit_math_h_l579_c3_8398_iffalse,
layer0_node51_MUX_bit_math_h_l579_c3_8398_return_output);

-- layer0_node52_MUX_bit_math_h_l590_c3_6d3d
layer0_node52_MUX_bit_math_h_l590_c3_6d3d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node52_MUX_bit_math_h_l590_c3_6d3d_cond,
layer0_node52_MUX_bit_math_h_l590_c3_6d3d_iftrue,
layer0_node52_MUX_bit_math_h_l590_c3_6d3d_iffalse,
layer0_node52_MUX_bit_math_h_l590_c3_6d3d_return_output);

-- layer0_node53_MUX_bit_math_h_l601_c3_6dc2
layer0_node53_MUX_bit_math_h_l601_c3_6dc2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node53_MUX_bit_math_h_l601_c3_6dc2_cond,
layer0_node53_MUX_bit_math_h_l601_c3_6dc2_iftrue,
layer0_node53_MUX_bit_math_h_l601_c3_6dc2_iffalse,
layer0_node53_MUX_bit_math_h_l601_c3_6dc2_return_output);

-- layer0_node54_MUX_bit_math_h_l612_c3_cab9
layer0_node54_MUX_bit_math_h_l612_c3_cab9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node54_MUX_bit_math_h_l612_c3_cab9_cond,
layer0_node54_MUX_bit_math_h_l612_c3_cab9_iftrue,
layer0_node54_MUX_bit_math_h_l612_c3_cab9_iffalse,
layer0_node54_MUX_bit_math_h_l612_c3_cab9_return_output);

-- layer0_node55_MUX_bit_math_h_l623_c3_2e5e
layer0_node55_MUX_bit_math_h_l623_c3_2e5e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node55_MUX_bit_math_h_l623_c3_2e5e_cond,
layer0_node55_MUX_bit_math_h_l623_c3_2e5e_iftrue,
layer0_node55_MUX_bit_math_h_l623_c3_2e5e_iffalse,
layer0_node55_MUX_bit_math_h_l623_c3_2e5e_return_output);

-- layer0_node56_MUX_bit_math_h_l634_c3_ab19
layer0_node56_MUX_bit_math_h_l634_c3_ab19 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node56_MUX_bit_math_h_l634_c3_ab19_cond,
layer0_node56_MUX_bit_math_h_l634_c3_ab19_iftrue,
layer0_node56_MUX_bit_math_h_l634_c3_ab19_iffalse,
layer0_node56_MUX_bit_math_h_l634_c3_ab19_return_output);

-- layer0_node57_MUX_bit_math_h_l645_c3_cec5
layer0_node57_MUX_bit_math_h_l645_c3_cec5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node57_MUX_bit_math_h_l645_c3_cec5_cond,
layer0_node57_MUX_bit_math_h_l645_c3_cec5_iftrue,
layer0_node57_MUX_bit_math_h_l645_c3_cec5_iffalse,
layer0_node57_MUX_bit_math_h_l645_c3_cec5_return_output);

-- layer0_node58_MUX_bit_math_h_l656_c3_312b
layer0_node58_MUX_bit_math_h_l656_c3_312b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node58_MUX_bit_math_h_l656_c3_312b_cond,
layer0_node58_MUX_bit_math_h_l656_c3_312b_iftrue,
layer0_node58_MUX_bit_math_h_l656_c3_312b_iffalse,
layer0_node58_MUX_bit_math_h_l656_c3_312b_return_output);

-- layer0_node59_MUX_bit_math_h_l667_c3_672d
layer0_node59_MUX_bit_math_h_l667_c3_672d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node59_MUX_bit_math_h_l667_c3_672d_cond,
layer0_node59_MUX_bit_math_h_l667_c3_672d_iftrue,
layer0_node59_MUX_bit_math_h_l667_c3_672d_iffalse,
layer0_node59_MUX_bit_math_h_l667_c3_672d_return_output);

-- layer0_node60_MUX_bit_math_h_l678_c3_9a42
layer0_node60_MUX_bit_math_h_l678_c3_9a42 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node60_MUX_bit_math_h_l678_c3_9a42_cond,
layer0_node60_MUX_bit_math_h_l678_c3_9a42_iftrue,
layer0_node60_MUX_bit_math_h_l678_c3_9a42_iffalse,
layer0_node60_MUX_bit_math_h_l678_c3_9a42_return_output);

-- layer0_node61_MUX_bit_math_h_l689_c3_be95
layer0_node61_MUX_bit_math_h_l689_c3_be95 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node61_MUX_bit_math_h_l689_c3_be95_cond,
layer0_node61_MUX_bit_math_h_l689_c3_be95_iftrue,
layer0_node61_MUX_bit_math_h_l689_c3_be95_iffalse,
layer0_node61_MUX_bit_math_h_l689_c3_be95_return_output);

-- layer0_node62_MUX_bit_math_h_l700_c3_8a98
layer0_node62_MUX_bit_math_h_l700_c3_8a98 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node62_MUX_bit_math_h_l700_c3_8a98_cond,
layer0_node62_MUX_bit_math_h_l700_c3_8a98_iftrue,
layer0_node62_MUX_bit_math_h_l700_c3_8a98_iffalse,
layer0_node62_MUX_bit_math_h_l700_c3_8a98_return_output);

-- layer0_node63_MUX_bit_math_h_l711_c3_45fc
layer0_node63_MUX_bit_math_h_l711_c3_45fc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node63_MUX_bit_math_h_l711_c3_45fc_cond,
layer0_node63_MUX_bit_math_h_l711_c3_45fc_iftrue,
layer0_node63_MUX_bit_math_h_l711_c3_45fc_iffalse,
layer0_node63_MUX_bit_math_h_l711_c3_45fc_return_output);

-- layer1_node0_MUX_bit_math_h_l728_c3_2ff0
layer1_node0_MUX_bit_math_h_l728_c3_2ff0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node0_MUX_bit_math_h_l728_c3_2ff0_cond,
layer1_node0_MUX_bit_math_h_l728_c3_2ff0_iftrue,
layer1_node0_MUX_bit_math_h_l728_c3_2ff0_iffalse,
layer1_node0_MUX_bit_math_h_l728_c3_2ff0_return_output);

-- layer1_node1_MUX_bit_math_h_l739_c3_8d8d
layer1_node1_MUX_bit_math_h_l739_c3_8d8d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node1_MUX_bit_math_h_l739_c3_8d8d_cond,
layer1_node1_MUX_bit_math_h_l739_c3_8d8d_iftrue,
layer1_node1_MUX_bit_math_h_l739_c3_8d8d_iffalse,
layer1_node1_MUX_bit_math_h_l739_c3_8d8d_return_output);

-- layer1_node2_MUX_bit_math_h_l750_c3_7ed6
layer1_node2_MUX_bit_math_h_l750_c3_7ed6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node2_MUX_bit_math_h_l750_c3_7ed6_cond,
layer1_node2_MUX_bit_math_h_l750_c3_7ed6_iftrue,
layer1_node2_MUX_bit_math_h_l750_c3_7ed6_iffalse,
layer1_node2_MUX_bit_math_h_l750_c3_7ed6_return_output);

-- layer1_node3_MUX_bit_math_h_l761_c3_68af
layer1_node3_MUX_bit_math_h_l761_c3_68af : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node3_MUX_bit_math_h_l761_c3_68af_cond,
layer1_node3_MUX_bit_math_h_l761_c3_68af_iftrue,
layer1_node3_MUX_bit_math_h_l761_c3_68af_iffalse,
layer1_node3_MUX_bit_math_h_l761_c3_68af_return_output);

-- layer1_node4_MUX_bit_math_h_l772_c3_e8c5
layer1_node4_MUX_bit_math_h_l772_c3_e8c5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node4_MUX_bit_math_h_l772_c3_e8c5_cond,
layer1_node4_MUX_bit_math_h_l772_c3_e8c5_iftrue,
layer1_node4_MUX_bit_math_h_l772_c3_e8c5_iffalse,
layer1_node4_MUX_bit_math_h_l772_c3_e8c5_return_output);

-- layer1_node5_MUX_bit_math_h_l783_c3_7ab9
layer1_node5_MUX_bit_math_h_l783_c3_7ab9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node5_MUX_bit_math_h_l783_c3_7ab9_cond,
layer1_node5_MUX_bit_math_h_l783_c3_7ab9_iftrue,
layer1_node5_MUX_bit_math_h_l783_c3_7ab9_iffalse,
layer1_node5_MUX_bit_math_h_l783_c3_7ab9_return_output);

-- layer1_node6_MUX_bit_math_h_l794_c3_1dbe
layer1_node6_MUX_bit_math_h_l794_c3_1dbe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node6_MUX_bit_math_h_l794_c3_1dbe_cond,
layer1_node6_MUX_bit_math_h_l794_c3_1dbe_iftrue,
layer1_node6_MUX_bit_math_h_l794_c3_1dbe_iffalse,
layer1_node6_MUX_bit_math_h_l794_c3_1dbe_return_output);

-- layer1_node7_MUX_bit_math_h_l805_c3_6dfe
layer1_node7_MUX_bit_math_h_l805_c3_6dfe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node7_MUX_bit_math_h_l805_c3_6dfe_cond,
layer1_node7_MUX_bit_math_h_l805_c3_6dfe_iftrue,
layer1_node7_MUX_bit_math_h_l805_c3_6dfe_iffalse,
layer1_node7_MUX_bit_math_h_l805_c3_6dfe_return_output);

-- layer1_node8_MUX_bit_math_h_l816_c3_5d19
layer1_node8_MUX_bit_math_h_l816_c3_5d19 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node8_MUX_bit_math_h_l816_c3_5d19_cond,
layer1_node8_MUX_bit_math_h_l816_c3_5d19_iftrue,
layer1_node8_MUX_bit_math_h_l816_c3_5d19_iffalse,
layer1_node8_MUX_bit_math_h_l816_c3_5d19_return_output);

-- layer1_node9_MUX_bit_math_h_l827_c3_fe3d
layer1_node9_MUX_bit_math_h_l827_c3_fe3d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node9_MUX_bit_math_h_l827_c3_fe3d_cond,
layer1_node9_MUX_bit_math_h_l827_c3_fe3d_iftrue,
layer1_node9_MUX_bit_math_h_l827_c3_fe3d_iffalse,
layer1_node9_MUX_bit_math_h_l827_c3_fe3d_return_output);

-- layer1_node10_MUX_bit_math_h_l838_c3_cc59
layer1_node10_MUX_bit_math_h_l838_c3_cc59 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node10_MUX_bit_math_h_l838_c3_cc59_cond,
layer1_node10_MUX_bit_math_h_l838_c3_cc59_iftrue,
layer1_node10_MUX_bit_math_h_l838_c3_cc59_iffalse,
layer1_node10_MUX_bit_math_h_l838_c3_cc59_return_output);

-- layer1_node11_MUX_bit_math_h_l849_c3_6ba8
layer1_node11_MUX_bit_math_h_l849_c3_6ba8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node11_MUX_bit_math_h_l849_c3_6ba8_cond,
layer1_node11_MUX_bit_math_h_l849_c3_6ba8_iftrue,
layer1_node11_MUX_bit_math_h_l849_c3_6ba8_iffalse,
layer1_node11_MUX_bit_math_h_l849_c3_6ba8_return_output);

-- layer1_node12_MUX_bit_math_h_l860_c3_e057
layer1_node12_MUX_bit_math_h_l860_c3_e057 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node12_MUX_bit_math_h_l860_c3_e057_cond,
layer1_node12_MUX_bit_math_h_l860_c3_e057_iftrue,
layer1_node12_MUX_bit_math_h_l860_c3_e057_iffalse,
layer1_node12_MUX_bit_math_h_l860_c3_e057_return_output);

-- layer1_node13_MUX_bit_math_h_l871_c3_aad3
layer1_node13_MUX_bit_math_h_l871_c3_aad3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node13_MUX_bit_math_h_l871_c3_aad3_cond,
layer1_node13_MUX_bit_math_h_l871_c3_aad3_iftrue,
layer1_node13_MUX_bit_math_h_l871_c3_aad3_iffalse,
layer1_node13_MUX_bit_math_h_l871_c3_aad3_return_output);

-- layer1_node14_MUX_bit_math_h_l882_c3_0d3c
layer1_node14_MUX_bit_math_h_l882_c3_0d3c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node14_MUX_bit_math_h_l882_c3_0d3c_cond,
layer1_node14_MUX_bit_math_h_l882_c3_0d3c_iftrue,
layer1_node14_MUX_bit_math_h_l882_c3_0d3c_iffalse,
layer1_node14_MUX_bit_math_h_l882_c3_0d3c_return_output);

-- layer1_node15_MUX_bit_math_h_l893_c3_6301
layer1_node15_MUX_bit_math_h_l893_c3_6301 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node15_MUX_bit_math_h_l893_c3_6301_cond,
layer1_node15_MUX_bit_math_h_l893_c3_6301_iftrue,
layer1_node15_MUX_bit_math_h_l893_c3_6301_iffalse,
layer1_node15_MUX_bit_math_h_l893_c3_6301_return_output);

-- layer1_node16_MUX_bit_math_h_l904_c3_60f0
layer1_node16_MUX_bit_math_h_l904_c3_60f0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node16_MUX_bit_math_h_l904_c3_60f0_cond,
layer1_node16_MUX_bit_math_h_l904_c3_60f0_iftrue,
layer1_node16_MUX_bit_math_h_l904_c3_60f0_iffalse,
layer1_node16_MUX_bit_math_h_l904_c3_60f0_return_output);

-- layer1_node17_MUX_bit_math_h_l915_c3_d47f
layer1_node17_MUX_bit_math_h_l915_c3_d47f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node17_MUX_bit_math_h_l915_c3_d47f_cond,
layer1_node17_MUX_bit_math_h_l915_c3_d47f_iftrue,
layer1_node17_MUX_bit_math_h_l915_c3_d47f_iffalse,
layer1_node17_MUX_bit_math_h_l915_c3_d47f_return_output);

-- layer1_node18_MUX_bit_math_h_l926_c3_678f
layer1_node18_MUX_bit_math_h_l926_c3_678f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node18_MUX_bit_math_h_l926_c3_678f_cond,
layer1_node18_MUX_bit_math_h_l926_c3_678f_iftrue,
layer1_node18_MUX_bit_math_h_l926_c3_678f_iffalse,
layer1_node18_MUX_bit_math_h_l926_c3_678f_return_output);

-- layer1_node19_MUX_bit_math_h_l937_c3_eb8f
layer1_node19_MUX_bit_math_h_l937_c3_eb8f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node19_MUX_bit_math_h_l937_c3_eb8f_cond,
layer1_node19_MUX_bit_math_h_l937_c3_eb8f_iftrue,
layer1_node19_MUX_bit_math_h_l937_c3_eb8f_iffalse,
layer1_node19_MUX_bit_math_h_l937_c3_eb8f_return_output);

-- layer1_node20_MUX_bit_math_h_l948_c3_588a
layer1_node20_MUX_bit_math_h_l948_c3_588a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node20_MUX_bit_math_h_l948_c3_588a_cond,
layer1_node20_MUX_bit_math_h_l948_c3_588a_iftrue,
layer1_node20_MUX_bit_math_h_l948_c3_588a_iffalse,
layer1_node20_MUX_bit_math_h_l948_c3_588a_return_output);

-- layer1_node21_MUX_bit_math_h_l959_c3_1823
layer1_node21_MUX_bit_math_h_l959_c3_1823 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node21_MUX_bit_math_h_l959_c3_1823_cond,
layer1_node21_MUX_bit_math_h_l959_c3_1823_iftrue,
layer1_node21_MUX_bit_math_h_l959_c3_1823_iffalse,
layer1_node21_MUX_bit_math_h_l959_c3_1823_return_output);

-- layer1_node22_MUX_bit_math_h_l970_c3_6904
layer1_node22_MUX_bit_math_h_l970_c3_6904 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node22_MUX_bit_math_h_l970_c3_6904_cond,
layer1_node22_MUX_bit_math_h_l970_c3_6904_iftrue,
layer1_node22_MUX_bit_math_h_l970_c3_6904_iffalse,
layer1_node22_MUX_bit_math_h_l970_c3_6904_return_output);

-- layer1_node23_MUX_bit_math_h_l981_c3_f890
layer1_node23_MUX_bit_math_h_l981_c3_f890 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node23_MUX_bit_math_h_l981_c3_f890_cond,
layer1_node23_MUX_bit_math_h_l981_c3_f890_iftrue,
layer1_node23_MUX_bit_math_h_l981_c3_f890_iffalse,
layer1_node23_MUX_bit_math_h_l981_c3_f890_return_output);

-- layer1_node24_MUX_bit_math_h_l992_c3_4e65
layer1_node24_MUX_bit_math_h_l992_c3_4e65 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node24_MUX_bit_math_h_l992_c3_4e65_cond,
layer1_node24_MUX_bit_math_h_l992_c3_4e65_iftrue,
layer1_node24_MUX_bit_math_h_l992_c3_4e65_iffalse,
layer1_node24_MUX_bit_math_h_l992_c3_4e65_return_output);

-- layer1_node25_MUX_bit_math_h_l1003_c3_f943
layer1_node25_MUX_bit_math_h_l1003_c3_f943 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node25_MUX_bit_math_h_l1003_c3_f943_cond,
layer1_node25_MUX_bit_math_h_l1003_c3_f943_iftrue,
layer1_node25_MUX_bit_math_h_l1003_c3_f943_iffalse,
layer1_node25_MUX_bit_math_h_l1003_c3_f943_return_output);

-- layer1_node26_MUX_bit_math_h_l1014_c3_aa20
layer1_node26_MUX_bit_math_h_l1014_c3_aa20 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node26_MUX_bit_math_h_l1014_c3_aa20_cond,
layer1_node26_MUX_bit_math_h_l1014_c3_aa20_iftrue,
layer1_node26_MUX_bit_math_h_l1014_c3_aa20_iffalse,
layer1_node26_MUX_bit_math_h_l1014_c3_aa20_return_output);

-- layer1_node27_MUX_bit_math_h_l1025_c3_a3a3
layer1_node27_MUX_bit_math_h_l1025_c3_a3a3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_cond,
layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_iftrue,
layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_iffalse,
layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_return_output);

-- layer1_node28_MUX_bit_math_h_l1036_c3_85a0
layer1_node28_MUX_bit_math_h_l1036_c3_85a0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node28_MUX_bit_math_h_l1036_c3_85a0_cond,
layer1_node28_MUX_bit_math_h_l1036_c3_85a0_iftrue,
layer1_node28_MUX_bit_math_h_l1036_c3_85a0_iffalse,
layer1_node28_MUX_bit_math_h_l1036_c3_85a0_return_output);

-- layer1_node29_MUX_bit_math_h_l1047_c3_953f
layer1_node29_MUX_bit_math_h_l1047_c3_953f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node29_MUX_bit_math_h_l1047_c3_953f_cond,
layer1_node29_MUX_bit_math_h_l1047_c3_953f_iftrue,
layer1_node29_MUX_bit_math_h_l1047_c3_953f_iffalse,
layer1_node29_MUX_bit_math_h_l1047_c3_953f_return_output);

-- layer1_node30_MUX_bit_math_h_l1058_c3_c3ba
layer1_node30_MUX_bit_math_h_l1058_c3_c3ba : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_cond,
layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_iftrue,
layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_iffalse,
layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_return_output);

-- layer1_node31_MUX_bit_math_h_l1069_c3_82fc
layer1_node31_MUX_bit_math_h_l1069_c3_82fc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node31_MUX_bit_math_h_l1069_c3_82fc_cond,
layer1_node31_MUX_bit_math_h_l1069_c3_82fc_iftrue,
layer1_node31_MUX_bit_math_h_l1069_c3_82fc_iffalse,
layer1_node31_MUX_bit_math_h_l1069_c3_82fc_return_output);

-- layer2_node0_MUX_bit_math_h_l1086_c3_4e60
layer2_node0_MUX_bit_math_h_l1086_c3_4e60 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node0_MUX_bit_math_h_l1086_c3_4e60_cond,
layer2_node0_MUX_bit_math_h_l1086_c3_4e60_iftrue,
layer2_node0_MUX_bit_math_h_l1086_c3_4e60_iffalse,
layer2_node0_MUX_bit_math_h_l1086_c3_4e60_return_output);

-- layer2_node1_MUX_bit_math_h_l1097_c3_12bb
layer2_node1_MUX_bit_math_h_l1097_c3_12bb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node1_MUX_bit_math_h_l1097_c3_12bb_cond,
layer2_node1_MUX_bit_math_h_l1097_c3_12bb_iftrue,
layer2_node1_MUX_bit_math_h_l1097_c3_12bb_iffalse,
layer2_node1_MUX_bit_math_h_l1097_c3_12bb_return_output);

-- layer2_node2_MUX_bit_math_h_l1108_c3_fcbb
layer2_node2_MUX_bit_math_h_l1108_c3_fcbb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_cond,
layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_iftrue,
layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_iffalse,
layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_return_output);

-- layer2_node3_MUX_bit_math_h_l1119_c3_8c7b
layer2_node3_MUX_bit_math_h_l1119_c3_8c7b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_cond,
layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_iftrue,
layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_iffalse,
layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_return_output);

-- layer2_node4_MUX_bit_math_h_l1130_c3_3de0
layer2_node4_MUX_bit_math_h_l1130_c3_3de0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node4_MUX_bit_math_h_l1130_c3_3de0_cond,
layer2_node4_MUX_bit_math_h_l1130_c3_3de0_iftrue,
layer2_node4_MUX_bit_math_h_l1130_c3_3de0_iffalse,
layer2_node4_MUX_bit_math_h_l1130_c3_3de0_return_output);

-- layer2_node5_MUX_bit_math_h_l1141_c3_a5f6
layer2_node5_MUX_bit_math_h_l1141_c3_a5f6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_cond,
layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_iftrue,
layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_iffalse,
layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_return_output);

-- layer2_node6_MUX_bit_math_h_l1152_c3_3828
layer2_node6_MUX_bit_math_h_l1152_c3_3828 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node6_MUX_bit_math_h_l1152_c3_3828_cond,
layer2_node6_MUX_bit_math_h_l1152_c3_3828_iftrue,
layer2_node6_MUX_bit_math_h_l1152_c3_3828_iffalse,
layer2_node6_MUX_bit_math_h_l1152_c3_3828_return_output);

-- layer2_node7_MUX_bit_math_h_l1163_c3_f226
layer2_node7_MUX_bit_math_h_l1163_c3_f226 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node7_MUX_bit_math_h_l1163_c3_f226_cond,
layer2_node7_MUX_bit_math_h_l1163_c3_f226_iftrue,
layer2_node7_MUX_bit_math_h_l1163_c3_f226_iffalse,
layer2_node7_MUX_bit_math_h_l1163_c3_f226_return_output);

-- layer2_node8_MUX_bit_math_h_l1174_c3_49b7
layer2_node8_MUX_bit_math_h_l1174_c3_49b7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node8_MUX_bit_math_h_l1174_c3_49b7_cond,
layer2_node8_MUX_bit_math_h_l1174_c3_49b7_iftrue,
layer2_node8_MUX_bit_math_h_l1174_c3_49b7_iffalse,
layer2_node8_MUX_bit_math_h_l1174_c3_49b7_return_output);

-- layer2_node9_MUX_bit_math_h_l1185_c3_934f
layer2_node9_MUX_bit_math_h_l1185_c3_934f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node9_MUX_bit_math_h_l1185_c3_934f_cond,
layer2_node9_MUX_bit_math_h_l1185_c3_934f_iftrue,
layer2_node9_MUX_bit_math_h_l1185_c3_934f_iffalse,
layer2_node9_MUX_bit_math_h_l1185_c3_934f_return_output);

-- layer2_node10_MUX_bit_math_h_l1196_c3_3f7c
layer2_node10_MUX_bit_math_h_l1196_c3_3f7c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_cond,
layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_iftrue,
layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_iffalse,
layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_return_output);

-- layer2_node11_MUX_bit_math_h_l1207_c3_d0a7
layer2_node11_MUX_bit_math_h_l1207_c3_d0a7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_cond,
layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_iftrue,
layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_iffalse,
layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_return_output);

-- layer2_node12_MUX_bit_math_h_l1218_c3_0726
layer2_node12_MUX_bit_math_h_l1218_c3_0726 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node12_MUX_bit_math_h_l1218_c3_0726_cond,
layer2_node12_MUX_bit_math_h_l1218_c3_0726_iftrue,
layer2_node12_MUX_bit_math_h_l1218_c3_0726_iffalse,
layer2_node12_MUX_bit_math_h_l1218_c3_0726_return_output);

-- layer2_node13_MUX_bit_math_h_l1229_c3_754d
layer2_node13_MUX_bit_math_h_l1229_c3_754d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node13_MUX_bit_math_h_l1229_c3_754d_cond,
layer2_node13_MUX_bit_math_h_l1229_c3_754d_iftrue,
layer2_node13_MUX_bit_math_h_l1229_c3_754d_iffalse,
layer2_node13_MUX_bit_math_h_l1229_c3_754d_return_output);

-- layer2_node14_MUX_bit_math_h_l1240_c3_2b9a
layer2_node14_MUX_bit_math_h_l1240_c3_2b9a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_cond,
layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_iftrue,
layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_iffalse,
layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_return_output);

-- layer2_node15_MUX_bit_math_h_l1251_c3_57b2
layer2_node15_MUX_bit_math_h_l1251_c3_57b2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node15_MUX_bit_math_h_l1251_c3_57b2_cond,
layer2_node15_MUX_bit_math_h_l1251_c3_57b2_iftrue,
layer2_node15_MUX_bit_math_h_l1251_c3_57b2_iffalse,
layer2_node15_MUX_bit_math_h_l1251_c3_57b2_return_output);

-- layer3_node0_MUX_bit_math_h_l1268_c3_e5cc
layer3_node0_MUX_bit_math_h_l1268_c3_e5cc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_cond,
layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_iftrue,
layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_iffalse,
layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_return_output);

-- layer3_node1_MUX_bit_math_h_l1279_c3_73ae
layer3_node1_MUX_bit_math_h_l1279_c3_73ae : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node1_MUX_bit_math_h_l1279_c3_73ae_cond,
layer3_node1_MUX_bit_math_h_l1279_c3_73ae_iftrue,
layer3_node1_MUX_bit_math_h_l1279_c3_73ae_iffalse,
layer3_node1_MUX_bit_math_h_l1279_c3_73ae_return_output);

-- layer3_node2_MUX_bit_math_h_l1290_c3_d8d2
layer3_node2_MUX_bit_math_h_l1290_c3_d8d2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_cond,
layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_iftrue,
layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_iffalse,
layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_return_output);

-- layer3_node3_MUX_bit_math_h_l1301_c3_827d
layer3_node3_MUX_bit_math_h_l1301_c3_827d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node3_MUX_bit_math_h_l1301_c3_827d_cond,
layer3_node3_MUX_bit_math_h_l1301_c3_827d_iftrue,
layer3_node3_MUX_bit_math_h_l1301_c3_827d_iffalse,
layer3_node3_MUX_bit_math_h_l1301_c3_827d_return_output);

-- layer3_node4_MUX_bit_math_h_l1312_c3_ca04
layer3_node4_MUX_bit_math_h_l1312_c3_ca04 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node4_MUX_bit_math_h_l1312_c3_ca04_cond,
layer3_node4_MUX_bit_math_h_l1312_c3_ca04_iftrue,
layer3_node4_MUX_bit_math_h_l1312_c3_ca04_iffalse,
layer3_node4_MUX_bit_math_h_l1312_c3_ca04_return_output);

-- layer3_node5_MUX_bit_math_h_l1323_c3_56dd
layer3_node5_MUX_bit_math_h_l1323_c3_56dd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node5_MUX_bit_math_h_l1323_c3_56dd_cond,
layer3_node5_MUX_bit_math_h_l1323_c3_56dd_iftrue,
layer3_node5_MUX_bit_math_h_l1323_c3_56dd_iffalse,
layer3_node5_MUX_bit_math_h_l1323_c3_56dd_return_output);

-- layer3_node6_MUX_bit_math_h_l1334_c3_07bd
layer3_node6_MUX_bit_math_h_l1334_c3_07bd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node6_MUX_bit_math_h_l1334_c3_07bd_cond,
layer3_node6_MUX_bit_math_h_l1334_c3_07bd_iftrue,
layer3_node6_MUX_bit_math_h_l1334_c3_07bd_iffalse,
layer3_node6_MUX_bit_math_h_l1334_c3_07bd_return_output);

-- layer3_node7_MUX_bit_math_h_l1345_c3_5a50
layer3_node7_MUX_bit_math_h_l1345_c3_5a50 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node7_MUX_bit_math_h_l1345_c3_5a50_cond,
layer3_node7_MUX_bit_math_h_l1345_c3_5a50_iftrue,
layer3_node7_MUX_bit_math_h_l1345_c3_5a50_iffalse,
layer3_node7_MUX_bit_math_h_l1345_c3_5a50_return_output);

-- layer4_node0_MUX_bit_math_h_l1362_c3_f5a3
layer4_node0_MUX_bit_math_h_l1362_c3_f5a3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_cond,
layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_iftrue,
layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_iffalse,
layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_return_output);

-- layer4_node1_MUX_bit_math_h_l1373_c3_402b
layer4_node1_MUX_bit_math_h_l1373_c3_402b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer4_node1_MUX_bit_math_h_l1373_c3_402b_cond,
layer4_node1_MUX_bit_math_h_l1373_c3_402b_iftrue,
layer4_node1_MUX_bit_math_h_l1373_c3_402b_iffalse,
layer4_node1_MUX_bit_math_h_l1373_c3_402b_return_output);

-- layer4_node2_MUX_bit_math_h_l1384_c3_5f80
layer4_node2_MUX_bit_math_h_l1384_c3_5f80 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer4_node2_MUX_bit_math_h_l1384_c3_5f80_cond,
layer4_node2_MUX_bit_math_h_l1384_c3_5f80_iftrue,
layer4_node2_MUX_bit_math_h_l1384_c3_5f80_iffalse,
layer4_node2_MUX_bit_math_h_l1384_c3_5f80_return_output);

-- layer4_node3_MUX_bit_math_h_l1395_c3_4d9c
layer4_node3_MUX_bit_math_h_l1395_c3_4d9c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_cond,
layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_iftrue,
layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_iffalse,
layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_return_output);

-- layer5_node0_MUX_bit_math_h_l1412_c3_19e3
layer5_node0_MUX_bit_math_h_l1412_c3_19e3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer5_node0_MUX_bit_math_h_l1412_c3_19e3_cond,
layer5_node0_MUX_bit_math_h_l1412_c3_19e3_iftrue,
layer5_node0_MUX_bit_math_h_l1412_c3_19e3_iffalse,
layer5_node0_MUX_bit_math_h_l1412_c3_19e3_return_output);

-- layer5_node1_MUX_bit_math_h_l1423_c3_11f1
layer5_node1_MUX_bit_math_h_l1423_c3_11f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer5_node1_MUX_bit_math_h_l1423_c3_11f1_cond,
layer5_node1_MUX_bit_math_h_l1423_c3_11f1_iftrue,
layer5_node1_MUX_bit_math_h_l1423_c3_11f1_iffalse,
layer5_node1_MUX_bit_math_h_l1423_c3_11f1_return_output);

-- layer6_node0_MUX_bit_math_h_l1440_c3_f906
layer6_node0_MUX_bit_math_h_l1440_c3_f906 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer6_node0_MUX_bit_math_h_l1440_c3_f906_cond,
layer6_node0_MUX_bit_math_h_l1440_c3_f906_iftrue,
layer6_node0_MUX_bit_math_h_l1440_c3_f906_iffalse,
layer6_node0_MUX_bit_math_h_l1440_c3_f906_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 sel,
 in0,
 in1,
 in2,
 in3,
 in4,
 in5,
 in6,
 in7,
 in8,
 in9,
 in10,
 in11,
 in12,
 in13,
 in14,
 in15,
 in16,
 in17,
 in18,
 in19,
 in20,
 in21,
 in22,
 in23,
 in24,
 in25,
 in26,
 in27,
 in28,
 in29,
 in30,
 in31,
 in32,
 in33,
 in34,
 in35,
 in36,
 in37,
 in38,
 in39,
 in40,
 in41,
 in42,
 in43,
 in44,
 in45,
 in46,
 in47,
 in48,
 in49,
 in50,
 in51,
 in52,
 in53,
 in54,
 in55,
 in56,
 in57,
 in58,
 in59,
 in60,
 in61,
 in62,
 in63,
 in64,
 in65,
 in66,
 in67,
 in68,
 in69,
 in70,
 in71,
 in72,
 in73,
 in74,
 in75,
 in76,
 in77,
 in78,
 in79,
 in80,
 in81,
 in82,
 in83,
 in84,
 in85,
 in86,
 in87,
 in88,
 in89,
 in90,
 in91,
 in92,
 in93,
 in94,
 in95,
 in96,
 in97,
 in98,
 in99,
 in100,
 in101,
 in102,
 in103,
 in104,
 in105,
 in106,
 in107,
 in108,
 in109,
 in110,
 in111,
 in112,
 in113,
 in114,
 in115,
 in116,
 in117,
 in118,
 in119,
 in120,
 in121,
 in122,
 in123,
 in124,
 in125,
 in126,
 in127,
 -- All submodule outputs
 layer0_node0_MUX_bit_math_h_l18_c3_5c06_return_output,
 layer0_node1_MUX_bit_math_h_l29_c3_fa46_return_output,
 layer0_node2_MUX_bit_math_h_l40_c3_f68a_return_output,
 layer0_node3_MUX_bit_math_h_l51_c3_b336_return_output,
 layer0_node4_MUX_bit_math_h_l62_c3_07e7_return_output,
 layer0_node5_MUX_bit_math_h_l73_c3_282b_return_output,
 layer0_node6_MUX_bit_math_h_l84_c3_62f1_return_output,
 layer0_node7_MUX_bit_math_h_l95_c3_567b_return_output,
 layer0_node8_MUX_bit_math_h_l106_c3_47e5_return_output,
 layer0_node9_MUX_bit_math_h_l117_c3_f097_return_output,
 layer0_node10_MUX_bit_math_h_l128_c3_0e6c_return_output,
 layer0_node11_MUX_bit_math_h_l139_c3_3ab9_return_output,
 layer0_node12_MUX_bit_math_h_l150_c3_e611_return_output,
 layer0_node13_MUX_bit_math_h_l161_c3_e037_return_output,
 layer0_node14_MUX_bit_math_h_l172_c3_ad25_return_output,
 layer0_node15_MUX_bit_math_h_l183_c3_dacd_return_output,
 layer0_node16_MUX_bit_math_h_l194_c3_5393_return_output,
 layer0_node17_MUX_bit_math_h_l205_c3_4246_return_output,
 layer0_node18_MUX_bit_math_h_l216_c3_2748_return_output,
 layer0_node19_MUX_bit_math_h_l227_c3_1dae_return_output,
 layer0_node20_MUX_bit_math_h_l238_c3_e7c7_return_output,
 layer0_node21_MUX_bit_math_h_l249_c3_8f8c_return_output,
 layer0_node22_MUX_bit_math_h_l260_c3_321e_return_output,
 layer0_node23_MUX_bit_math_h_l271_c3_86c3_return_output,
 layer0_node24_MUX_bit_math_h_l282_c3_2992_return_output,
 layer0_node25_MUX_bit_math_h_l293_c3_ece2_return_output,
 layer0_node26_MUX_bit_math_h_l304_c3_7f9b_return_output,
 layer0_node27_MUX_bit_math_h_l315_c3_5c0f_return_output,
 layer0_node28_MUX_bit_math_h_l326_c3_12a3_return_output,
 layer0_node29_MUX_bit_math_h_l337_c3_cbb8_return_output,
 layer0_node30_MUX_bit_math_h_l348_c3_8c5c_return_output,
 layer0_node31_MUX_bit_math_h_l359_c3_d6b9_return_output,
 layer0_node32_MUX_bit_math_h_l370_c3_3d24_return_output,
 layer0_node33_MUX_bit_math_h_l381_c3_bdd0_return_output,
 layer0_node34_MUX_bit_math_h_l392_c3_f617_return_output,
 layer0_node35_MUX_bit_math_h_l403_c3_683e_return_output,
 layer0_node36_MUX_bit_math_h_l414_c3_cd2c_return_output,
 layer0_node37_MUX_bit_math_h_l425_c3_2485_return_output,
 layer0_node38_MUX_bit_math_h_l436_c3_c940_return_output,
 layer0_node39_MUX_bit_math_h_l447_c3_b150_return_output,
 layer0_node40_MUX_bit_math_h_l458_c3_c977_return_output,
 layer0_node41_MUX_bit_math_h_l469_c3_b3bf_return_output,
 layer0_node42_MUX_bit_math_h_l480_c3_c677_return_output,
 layer0_node43_MUX_bit_math_h_l491_c3_2838_return_output,
 layer0_node44_MUX_bit_math_h_l502_c3_6b96_return_output,
 layer0_node45_MUX_bit_math_h_l513_c3_b86e_return_output,
 layer0_node46_MUX_bit_math_h_l524_c3_4ef5_return_output,
 layer0_node47_MUX_bit_math_h_l535_c3_21f3_return_output,
 layer0_node48_MUX_bit_math_h_l546_c3_5be4_return_output,
 layer0_node49_MUX_bit_math_h_l557_c3_3410_return_output,
 layer0_node50_MUX_bit_math_h_l568_c3_4522_return_output,
 layer0_node51_MUX_bit_math_h_l579_c3_8398_return_output,
 layer0_node52_MUX_bit_math_h_l590_c3_6d3d_return_output,
 layer0_node53_MUX_bit_math_h_l601_c3_6dc2_return_output,
 layer0_node54_MUX_bit_math_h_l612_c3_cab9_return_output,
 layer0_node55_MUX_bit_math_h_l623_c3_2e5e_return_output,
 layer0_node56_MUX_bit_math_h_l634_c3_ab19_return_output,
 layer0_node57_MUX_bit_math_h_l645_c3_cec5_return_output,
 layer0_node58_MUX_bit_math_h_l656_c3_312b_return_output,
 layer0_node59_MUX_bit_math_h_l667_c3_672d_return_output,
 layer0_node60_MUX_bit_math_h_l678_c3_9a42_return_output,
 layer0_node61_MUX_bit_math_h_l689_c3_be95_return_output,
 layer0_node62_MUX_bit_math_h_l700_c3_8a98_return_output,
 layer0_node63_MUX_bit_math_h_l711_c3_45fc_return_output,
 layer1_node0_MUX_bit_math_h_l728_c3_2ff0_return_output,
 layer1_node1_MUX_bit_math_h_l739_c3_8d8d_return_output,
 layer1_node2_MUX_bit_math_h_l750_c3_7ed6_return_output,
 layer1_node3_MUX_bit_math_h_l761_c3_68af_return_output,
 layer1_node4_MUX_bit_math_h_l772_c3_e8c5_return_output,
 layer1_node5_MUX_bit_math_h_l783_c3_7ab9_return_output,
 layer1_node6_MUX_bit_math_h_l794_c3_1dbe_return_output,
 layer1_node7_MUX_bit_math_h_l805_c3_6dfe_return_output,
 layer1_node8_MUX_bit_math_h_l816_c3_5d19_return_output,
 layer1_node9_MUX_bit_math_h_l827_c3_fe3d_return_output,
 layer1_node10_MUX_bit_math_h_l838_c3_cc59_return_output,
 layer1_node11_MUX_bit_math_h_l849_c3_6ba8_return_output,
 layer1_node12_MUX_bit_math_h_l860_c3_e057_return_output,
 layer1_node13_MUX_bit_math_h_l871_c3_aad3_return_output,
 layer1_node14_MUX_bit_math_h_l882_c3_0d3c_return_output,
 layer1_node15_MUX_bit_math_h_l893_c3_6301_return_output,
 layer1_node16_MUX_bit_math_h_l904_c3_60f0_return_output,
 layer1_node17_MUX_bit_math_h_l915_c3_d47f_return_output,
 layer1_node18_MUX_bit_math_h_l926_c3_678f_return_output,
 layer1_node19_MUX_bit_math_h_l937_c3_eb8f_return_output,
 layer1_node20_MUX_bit_math_h_l948_c3_588a_return_output,
 layer1_node21_MUX_bit_math_h_l959_c3_1823_return_output,
 layer1_node22_MUX_bit_math_h_l970_c3_6904_return_output,
 layer1_node23_MUX_bit_math_h_l981_c3_f890_return_output,
 layer1_node24_MUX_bit_math_h_l992_c3_4e65_return_output,
 layer1_node25_MUX_bit_math_h_l1003_c3_f943_return_output,
 layer1_node26_MUX_bit_math_h_l1014_c3_aa20_return_output,
 layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_return_output,
 layer1_node28_MUX_bit_math_h_l1036_c3_85a0_return_output,
 layer1_node29_MUX_bit_math_h_l1047_c3_953f_return_output,
 layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_return_output,
 layer1_node31_MUX_bit_math_h_l1069_c3_82fc_return_output,
 layer2_node0_MUX_bit_math_h_l1086_c3_4e60_return_output,
 layer2_node1_MUX_bit_math_h_l1097_c3_12bb_return_output,
 layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_return_output,
 layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_return_output,
 layer2_node4_MUX_bit_math_h_l1130_c3_3de0_return_output,
 layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_return_output,
 layer2_node6_MUX_bit_math_h_l1152_c3_3828_return_output,
 layer2_node7_MUX_bit_math_h_l1163_c3_f226_return_output,
 layer2_node8_MUX_bit_math_h_l1174_c3_49b7_return_output,
 layer2_node9_MUX_bit_math_h_l1185_c3_934f_return_output,
 layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_return_output,
 layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_return_output,
 layer2_node12_MUX_bit_math_h_l1218_c3_0726_return_output,
 layer2_node13_MUX_bit_math_h_l1229_c3_754d_return_output,
 layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_return_output,
 layer2_node15_MUX_bit_math_h_l1251_c3_57b2_return_output,
 layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_return_output,
 layer3_node1_MUX_bit_math_h_l1279_c3_73ae_return_output,
 layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_return_output,
 layer3_node3_MUX_bit_math_h_l1301_c3_827d_return_output,
 layer3_node4_MUX_bit_math_h_l1312_c3_ca04_return_output,
 layer3_node5_MUX_bit_math_h_l1323_c3_56dd_return_output,
 layer3_node6_MUX_bit_math_h_l1334_c3_07bd_return_output,
 layer3_node7_MUX_bit_math_h_l1345_c3_5a50_return_output,
 layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_return_output,
 layer4_node1_MUX_bit_math_h_l1373_c3_402b_return_output,
 layer4_node2_MUX_bit_math_h_l1384_c3_5f80_return_output,
 layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_return_output,
 layer5_node0_MUX_bit_math_h_l1412_c3_19e3_return_output,
 layer5_node1_MUX_bit_math_h_l1423_c3_11f1_return_output,
 layer6_node0_MUX_bit_math_h_l1440_c3_f906_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(7 downto 0);
 variable VAR_sel : unsigned(6 downto 0);
 variable VAR_in0 : unsigned(7 downto 0);
 variable VAR_in1 : unsigned(7 downto 0);
 variable VAR_in2 : unsigned(7 downto 0);
 variable VAR_in3 : unsigned(7 downto 0);
 variable VAR_in4 : unsigned(7 downto 0);
 variable VAR_in5 : unsigned(7 downto 0);
 variable VAR_in6 : unsigned(7 downto 0);
 variable VAR_in7 : unsigned(7 downto 0);
 variable VAR_in8 : unsigned(7 downto 0);
 variable VAR_in9 : unsigned(7 downto 0);
 variable VAR_in10 : unsigned(7 downto 0);
 variable VAR_in11 : unsigned(7 downto 0);
 variable VAR_in12 : unsigned(7 downto 0);
 variable VAR_in13 : unsigned(7 downto 0);
 variable VAR_in14 : unsigned(7 downto 0);
 variable VAR_in15 : unsigned(7 downto 0);
 variable VAR_in16 : unsigned(7 downto 0);
 variable VAR_in17 : unsigned(7 downto 0);
 variable VAR_in18 : unsigned(7 downto 0);
 variable VAR_in19 : unsigned(7 downto 0);
 variable VAR_in20 : unsigned(7 downto 0);
 variable VAR_in21 : unsigned(7 downto 0);
 variable VAR_in22 : unsigned(7 downto 0);
 variable VAR_in23 : unsigned(7 downto 0);
 variable VAR_in24 : unsigned(7 downto 0);
 variable VAR_in25 : unsigned(7 downto 0);
 variable VAR_in26 : unsigned(7 downto 0);
 variable VAR_in27 : unsigned(7 downto 0);
 variable VAR_in28 : unsigned(7 downto 0);
 variable VAR_in29 : unsigned(7 downto 0);
 variable VAR_in30 : unsigned(7 downto 0);
 variable VAR_in31 : unsigned(7 downto 0);
 variable VAR_in32 : unsigned(7 downto 0);
 variable VAR_in33 : unsigned(7 downto 0);
 variable VAR_in34 : unsigned(7 downto 0);
 variable VAR_in35 : unsigned(7 downto 0);
 variable VAR_in36 : unsigned(7 downto 0);
 variable VAR_in37 : unsigned(7 downto 0);
 variable VAR_in38 : unsigned(7 downto 0);
 variable VAR_in39 : unsigned(7 downto 0);
 variable VAR_in40 : unsigned(7 downto 0);
 variable VAR_in41 : unsigned(7 downto 0);
 variable VAR_in42 : unsigned(7 downto 0);
 variable VAR_in43 : unsigned(7 downto 0);
 variable VAR_in44 : unsigned(7 downto 0);
 variable VAR_in45 : unsigned(7 downto 0);
 variable VAR_in46 : unsigned(7 downto 0);
 variable VAR_in47 : unsigned(7 downto 0);
 variable VAR_in48 : unsigned(7 downto 0);
 variable VAR_in49 : unsigned(7 downto 0);
 variable VAR_in50 : unsigned(7 downto 0);
 variable VAR_in51 : unsigned(7 downto 0);
 variable VAR_in52 : unsigned(7 downto 0);
 variable VAR_in53 : unsigned(7 downto 0);
 variable VAR_in54 : unsigned(7 downto 0);
 variable VAR_in55 : unsigned(7 downto 0);
 variable VAR_in56 : unsigned(7 downto 0);
 variable VAR_in57 : unsigned(7 downto 0);
 variable VAR_in58 : unsigned(7 downto 0);
 variable VAR_in59 : unsigned(7 downto 0);
 variable VAR_in60 : unsigned(7 downto 0);
 variable VAR_in61 : unsigned(7 downto 0);
 variable VAR_in62 : unsigned(7 downto 0);
 variable VAR_in63 : unsigned(7 downto 0);
 variable VAR_in64 : unsigned(7 downto 0);
 variable VAR_in65 : unsigned(7 downto 0);
 variable VAR_in66 : unsigned(7 downto 0);
 variable VAR_in67 : unsigned(7 downto 0);
 variable VAR_in68 : unsigned(7 downto 0);
 variable VAR_in69 : unsigned(7 downto 0);
 variable VAR_in70 : unsigned(7 downto 0);
 variable VAR_in71 : unsigned(7 downto 0);
 variable VAR_in72 : unsigned(7 downto 0);
 variable VAR_in73 : unsigned(7 downto 0);
 variable VAR_in74 : unsigned(7 downto 0);
 variable VAR_in75 : unsigned(7 downto 0);
 variable VAR_in76 : unsigned(7 downto 0);
 variable VAR_in77 : unsigned(7 downto 0);
 variable VAR_in78 : unsigned(7 downto 0);
 variable VAR_in79 : unsigned(7 downto 0);
 variable VAR_in80 : unsigned(7 downto 0);
 variable VAR_in81 : unsigned(7 downto 0);
 variable VAR_in82 : unsigned(7 downto 0);
 variable VAR_in83 : unsigned(7 downto 0);
 variable VAR_in84 : unsigned(7 downto 0);
 variable VAR_in85 : unsigned(7 downto 0);
 variable VAR_in86 : unsigned(7 downto 0);
 variable VAR_in87 : unsigned(7 downto 0);
 variable VAR_in88 : unsigned(7 downto 0);
 variable VAR_in89 : unsigned(7 downto 0);
 variable VAR_in90 : unsigned(7 downto 0);
 variable VAR_in91 : unsigned(7 downto 0);
 variable VAR_in92 : unsigned(7 downto 0);
 variable VAR_in93 : unsigned(7 downto 0);
 variable VAR_in94 : unsigned(7 downto 0);
 variable VAR_in95 : unsigned(7 downto 0);
 variable VAR_in96 : unsigned(7 downto 0);
 variable VAR_in97 : unsigned(7 downto 0);
 variable VAR_in98 : unsigned(7 downto 0);
 variable VAR_in99 : unsigned(7 downto 0);
 variable VAR_in100 : unsigned(7 downto 0);
 variable VAR_in101 : unsigned(7 downto 0);
 variable VAR_in102 : unsigned(7 downto 0);
 variable VAR_in103 : unsigned(7 downto 0);
 variable VAR_in104 : unsigned(7 downto 0);
 variable VAR_in105 : unsigned(7 downto 0);
 variable VAR_in106 : unsigned(7 downto 0);
 variable VAR_in107 : unsigned(7 downto 0);
 variable VAR_in108 : unsigned(7 downto 0);
 variable VAR_in109 : unsigned(7 downto 0);
 variable VAR_in110 : unsigned(7 downto 0);
 variable VAR_in111 : unsigned(7 downto 0);
 variable VAR_in112 : unsigned(7 downto 0);
 variable VAR_in113 : unsigned(7 downto 0);
 variable VAR_in114 : unsigned(7 downto 0);
 variable VAR_in115 : unsigned(7 downto 0);
 variable VAR_in116 : unsigned(7 downto 0);
 variable VAR_in117 : unsigned(7 downto 0);
 variable VAR_in118 : unsigned(7 downto 0);
 variable VAR_in119 : unsigned(7 downto 0);
 variable VAR_in120 : unsigned(7 downto 0);
 variable VAR_in121 : unsigned(7 downto 0);
 variable VAR_in122 : unsigned(7 downto 0);
 variable VAR_in123 : unsigned(7 downto 0);
 variable VAR_in124 : unsigned(7 downto 0);
 variable VAR_in125 : unsigned(7 downto 0);
 variable VAR_in126 : unsigned(7 downto 0);
 variable VAR_in127 : unsigned(7 downto 0);
 variable VAR_sel0 : unsigned(0 downto 0);
 variable VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output : unsigned(0 downto 0);
 variable VAR_layer0_node0 : unsigned(7 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_5c06_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_5c06_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_5c06_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_5c06_cond : unsigned(0 downto 0);
 variable VAR_layer0_node1 : unsigned(7 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_fa46_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_fa46_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_fa46_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_fa46_cond : unsigned(0 downto 0);
 variable VAR_layer0_node2 : unsigned(7 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_f68a_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_f68a_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_f68a_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_f68a_cond : unsigned(0 downto 0);
 variable VAR_layer0_node3 : unsigned(7 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_b336_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_b336_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_b336_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_b336_cond : unsigned(0 downto 0);
 variable VAR_layer0_node4 : unsigned(7 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_07e7_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_07e7_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_07e7_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_07e7_cond : unsigned(0 downto 0);
 variable VAR_layer0_node5 : unsigned(7 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_282b_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_282b_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_282b_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_282b_cond : unsigned(0 downto 0);
 variable VAR_layer0_node6 : unsigned(7 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_62f1_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_62f1_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_62f1_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_62f1_cond : unsigned(0 downto 0);
 variable VAR_layer0_node7 : unsigned(7 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_567b_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_567b_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_567b_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_567b_cond : unsigned(0 downto 0);
 variable VAR_layer0_node8 : unsigned(7 downto 0);
 variable VAR_layer0_node8_MUX_bit_math_h_l106_c3_47e5_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node8_MUX_bit_math_h_l106_c3_47e5_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node8_MUX_bit_math_h_l106_c3_47e5_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node8_MUX_bit_math_h_l106_c3_47e5_cond : unsigned(0 downto 0);
 variable VAR_layer0_node9 : unsigned(7 downto 0);
 variable VAR_layer0_node9_MUX_bit_math_h_l117_c3_f097_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node9_MUX_bit_math_h_l117_c3_f097_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node9_MUX_bit_math_h_l117_c3_f097_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node9_MUX_bit_math_h_l117_c3_f097_cond : unsigned(0 downto 0);
 variable VAR_layer0_node10 : unsigned(7 downto 0);
 variable VAR_layer0_node10_MUX_bit_math_h_l128_c3_0e6c_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node10_MUX_bit_math_h_l128_c3_0e6c_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node10_MUX_bit_math_h_l128_c3_0e6c_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node10_MUX_bit_math_h_l128_c3_0e6c_cond : unsigned(0 downto 0);
 variable VAR_layer0_node11 : unsigned(7 downto 0);
 variable VAR_layer0_node11_MUX_bit_math_h_l139_c3_3ab9_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node11_MUX_bit_math_h_l139_c3_3ab9_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node11_MUX_bit_math_h_l139_c3_3ab9_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node11_MUX_bit_math_h_l139_c3_3ab9_cond : unsigned(0 downto 0);
 variable VAR_layer0_node12 : unsigned(7 downto 0);
 variable VAR_layer0_node12_MUX_bit_math_h_l150_c3_e611_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node12_MUX_bit_math_h_l150_c3_e611_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node12_MUX_bit_math_h_l150_c3_e611_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node12_MUX_bit_math_h_l150_c3_e611_cond : unsigned(0 downto 0);
 variable VAR_layer0_node13 : unsigned(7 downto 0);
 variable VAR_layer0_node13_MUX_bit_math_h_l161_c3_e037_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node13_MUX_bit_math_h_l161_c3_e037_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node13_MUX_bit_math_h_l161_c3_e037_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node13_MUX_bit_math_h_l161_c3_e037_cond : unsigned(0 downto 0);
 variable VAR_layer0_node14 : unsigned(7 downto 0);
 variable VAR_layer0_node14_MUX_bit_math_h_l172_c3_ad25_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node14_MUX_bit_math_h_l172_c3_ad25_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node14_MUX_bit_math_h_l172_c3_ad25_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node14_MUX_bit_math_h_l172_c3_ad25_cond : unsigned(0 downto 0);
 variable VAR_layer0_node15 : unsigned(7 downto 0);
 variable VAR_layer0_node15_MUX_bit_math_h_l183_c3_dacd_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node15_MUX_bit_math_h_l183_c3_dacd_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node15_MUX_bit_math_h_l183_c3_dacd_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node15_MUX_bit_math_h_l183_c3_dacd_cond : unsigned(0 downto 0);
 variable VAR_layer0_node16 : unsigned(7 downto 0);
 variable VAR_layer0_node16_MUX_bit_math_h_l194_c3_5393_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node16_MUX_bit_math_h_l194_c3_5393_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node16_MUX_bit_math_h_l194_c3_5393_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node16_MUX_bit_math_h_l194_c3_5393_cond : unsigned(0 downto 0);
 variable VAR_layer0_node17 : unsigned(7 downto 0);
 variable VAR_layer0_node17_MUX_bit_math_h_l205_c3_4246_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node17_MUX_bit_math_h_l205_c3_4246_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node17_MUX_bit_math_h_l205_c3_4246_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node17_MUX_bit_math_h_l205_c3_4246_cond : unsigned(0 downto 0);
 variable VAR_layer0_node18 : unsigned(7 downto 0);
 variable VAR_layer0_node18_MUX_bit_math_h_l216_c3_2748_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node18_MUX_bit_math_h_l216_c3_2748_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node18_MUX_bit_math_h_l216_c3_2748_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node18_MUX_bit_math_h_l216_c3_2748_cond : unsigned(0 downto 0);
 variable VAR_layer0_node19 : unsigned(7 downto 0);
 variable VAR_layer0_node19_MUX_bit_math_h_l227_c3_1dae_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node19_MUX_bit_math_h_l227_c3_1dae_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node19_MUX_bit_math_h_l227_c3_1dae_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node19_MUX_bit_math_h_l227_c3_1dae_cond : unsigned(0 downto 0);
 variable VAR_layer0_node20 : unsigned(7 downto 0);
 variable VAR_layer0_node20_MUX_bit_math_h_l238_c3_e7c7_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node20_MUX_bit_math_h_l238_c3_e7c7_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node20_MUX_bit_math_h_l238_c3_e7c7_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node20_MUX_bit_math_h_l238_c3_e7c7_cond : unsigned(0 downto 0);
 variable VAR_layer0_node21 : unsigned(7 downto 0);
 variable VAR_layer0_node21_MUX_bit_math_h_l249_c3_8f8c_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node21_MUX_bit_math_h_l249_c3_8f8c_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node21_MUX_bit_math_h_l249_c3_8f8c_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node21_MUX_bit_math_h_l249_c3_8f8c_cond : unsigned(0 downto 0);
 variable VAR_layer0_node22 : unsigned(7 downto 0);
 variable VAR_layer0_node22_MUX_bit_math_h_l260_c3_321e_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node22_MUX_bit_math_h_l260_c3_321e_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node22_MUX_bit_math_h_l260_c3_321e_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node22_MUX_bit_math_h_l260_c3_321e_cond : unsigned(0 downto 0);
 variable VAR_layer0_node23 : unsigned(7 downto 0);
 variable VAR_layer0_node23_MUX_bit_math_h_l271_c3_86c3_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node23_MUX_bit_math_h_l271_c3_86c3_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node23_MUX_bit_math_h_l271_c3_86c3_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node23_MUX_bit_math_h_l271_c3_86c3_cond : unsigned(0 downto 0);
 variable VAR_layer0_node24 : unsigned(7 downto 0);
 variable VAR_layer0_node24_MUX_bit_math_h_l282_c3_2992_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node24_MUX_bit_math_h_l282_c3_2992_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node24_MUX_bit_math_h_l282_c3_2992_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node24_MUX_bit_math_h_l282_c3_2992_cond : unsigned(0 downto 0);
 variable VAR_layer0_node25 : unsigned(7 downto 0);
 variable VAR_layer0_node25_MUX_bit_math_h_l293_c3_ece2_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node25_MUX_bit_math_h_l293_c3_ece2_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node25_MUX_bit_math_h_l293_c3_ece2_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node25_MUX_bit_math_h_l293_c3_ece2_cond : unsigned(0 downto 0);
 variable VAR_layer0_node26 : unsigned(7 downto 0);
 variable VAR_layer0_node26_MUX_bit_math_h_l304_c3_7f9b_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node26_MUX_bit_math_h_l304_c3_7f9b_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node26_MUX_bit_math_h_l304_c3_7f9b_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node26_MUX_bit_math_h_l304_c3_7f9b_cond : unsigned(0 downto 0);
 variable VAR_layer0_node27 : unsigned(7 downto 0);
 variable VAR_layer0_node27_MUX_bit_math_h_l315_c3_5c0f_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node27_MUX_bit_math_h_l315_c3_5c0f_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node27_MUX_bit_math_h_l315_c3_5c0f_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node27_MUX_bit_math_h_l315_c3_5c0f_cond : unsigned(0 downto 0);
 variable VAR_layer0_node28 : unsigned(7 downto 0);
 variable VAR_layer0_node28_MUX_bit_math_h_l326_c3_12a3_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node28_MUX_bit_math_h_l326_c3_12a3_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node28_MUX_bit_math_h_l326_c3_12a3_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node28_MUX_bit_math_h_l326_c3_12a3_cond : unsigned(0 downto 0);
 variable VAR_layer0_node29 : unsigned(7 downto 0);
 variable VAR_layer0_node29_MUX_bit_math_h_l337_c3_cbb8_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node29_MUX_bit_math_h_l337_c3_cbb8_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node29_MUX_bit_math_h_l337_c3_cbb8_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node29_MUX_bit_math_h_l337_c3_cbb8_cond : unsigned(0 downto 0);
 variable VAR_layer0_node30 : unsigned(7 downto 0);
 variable VAR_layer0_node30_MUX_bit_math_h_l348_c3_8c5c_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node30_MUX_bit_math_h_l348_c3_8c5c_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node30_MUX_bit_math_h_l348_c3_8c5c_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node30_MUX_bit_math_h_l348_c3_8c5c_cond : unsigned(0 downto 0);
 variable VAR_layer0_node31 : unsigned(7 downto 0);
 variable VAR_layer0_node31_MUX_bit_math_h_l359_c3_d6b9_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node31_MUX_bit_math_h_l359_c3_d6b9_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node31_MUX_bit_math_h_l359_c3_d6b9_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node31_MUX_bit_math_h_l359_c3_d6b9_cond : unsigned(0 downto 0);
 variable VAR_layer0_node32 : unsigned(7 downto 0);
 variable VAR_layer0_node32_MUX_bit_math_h_l370_c3_3d24_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node32_MUX_bit_math_h_l370_c3_3d24_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node32_MUX_bit_math_h_l370_c3_3d24_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node32_MUX_bit_math_h_l370_c3_3d24_cond : unsigned(0 downto 0);
 variable VAR_layer0_node33 : unsigned(7 downto 0);
 variable VAR_layer0_node33_MUX_bit_math_h_l381_c3_bdd0_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node33_MUX_bit_math_h_l381_c3_bdd0_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node33_MUX_bit_math_h_l381_c3_bdd0_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node33_MUX_bit_math_h_l381_c3_bdd0_cond : unsigned(0 downto 0);
 variable VAR_layer0_node34 : unsigned(7 downto 0);
 variable VAR_layer0_node34_MUX_bit_math_h_l392_c3_f617_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node34_MUX_bit_math_h_l392_c3_f617_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node34_MUX_bit_math_h_l392_c3_f617_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node34_MUX_bit_math_h_l392_c3_f617_cond : unsigned(0 downto 0);
 variable VAR_layer0_node35 : unsigned(7 downto 0);
 variable VAR_layer0_node35_MUX_bit_math_h_l403_c3_683e_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node35_MUX_bit_math_h_l403_c3_683e_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node35_MUX_bit_math_h_l403_c3_683e_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node35_MUX_bit_math_h_l403_c3_683e_cond : unsigned(0 downto 0);
 variable VAR_layer0_node36 : unsigned(7 downto 0);
 variable VAR_layer0_node36_MUX_bit_math_h_l414_c3_cd2c_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node36_MUX_bit_math_h_l414_c3_cd2c_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node36_MUX_bit_math_h_l414_c3_cd2c_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node36_MUX_bit_math_h_l414_c3_cd2c_cond : unsigned(0 downto 0);
 variable VAR_layer0_node37 : unsigned(7 downto 0);
 variable VAR_layer0_node37_MUX_bit_math_h_l425_c3_2485_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node37_MUX_bit_math_h_l425_c3_2485_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node37_MUX_bit_math_h_l425_c3_2485_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node37_MUX_bit_math_h_l425_c3_2485_cond : unsigned(0 downto 0);
 variable VAR_layer0_node38 : unsigned(7 downto 0);
 variable VAR_layer0_node38_MUX_bit_math_h_l436_c3_c940_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node38_MUX_bit_math_h_l436_c3_c940_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node38_MUX_bit_math_h_l436_c3_c940_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node38_MUX_bit_math_h_l436_c3_c940_cond : unsigned(0 downto 0);
 variable VAR_layer0_node39 : unsigned(7 downto 0);
 variable VAR_layer0_node39_MUX_bit_math_h_l447_c3_b150_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node39_MUX_bit_math_h_l447_c3_b150_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node39_MUX_bit_math_h_l447_c3_b150_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node39_MUX_bit_math_h_l447_c3_b150_cond : unsigned(0 downto 0);
 variable VAR_layer0_node40 : unsigned(7 downto 0);
 variable VAR_layer0_node40_MUX_bit_math_h_l458_c3_c977_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node40_MUX_bit_math_h_l458_c3_c977_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node40_MUX_bit_math_h_l458_c3_c977_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node40_MUX_bit_math_h_l458_c3_c977_cond : unsigned(0 downto 0);
 variable VAR_layer0_node41 : unsigned(7 downto 0);
 variable VAR_layer0_node41_MUX_bit_math_h_l469_c3_b3bf_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node41_MUX_bit_math_h_l469_c3_b3bf_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node41_MUX_bit_math_h_l469_c3_b3bf_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node41_MUX_bit_math_h_l469_c3_b3bf_cond : unsigned(0 downto 0);
 variable VAR_layer0_node42 : unsigned(7 downto 0);
 variable VAR_layer0_node42_MUX_bit_math_h_l480_c3_c677_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node42_MUX_bit_math_h_l480_c3_c677_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node42_MUX_bit_math_h_l480_c3_c677_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node42_MUX_bit_math_h_l480_c3_c677_cond : unsigned(0 downto 0);
 variable VAR_layer0_node43 : unsigned(7 downto 0);
 variable VAR_layer0_node43_MUX_bit_math_h_l491_c3_2838_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node43_MUX_bit_math_h_l491_c3_2838_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node43_MUX_bit_math_h_l491_c3_2838_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node43_MUX_bit_math_h_l491_c3_2838_cond : unsigned(0 downto 0);
 variable VAR_layer0_node44 : unsigned(7 downto 0);
 variable VAR_layer0_node44_MUX_bit_math_h_l502_c3_6b96_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node44_MUX_bit_math_h_l502_c3_6b96_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node44_MUX_bit_math_h_l502_c3_6b96_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node44_MUX_bit_math_h_l502_c3_6b96_cond : unsigned(0 downto 0);
 variable VAR_layer0_node45 : unsigned(7 downto 0);
 variable VAR_layer0_node45_MUX_bit_math_h_l513_c3_b86e_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node45_MUX_bit_math_h_l513_c3_b86e_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node45_MUX_bit_math_h_l513_c3_b86e_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node45_MUX_bit_math_h_l513_c3_b86e_cond : unsigned(0 downto 0);
 variable VAR_layer0_node46 : unsigned(7 downto 0);
 variable VAR_layer0_node46_MUX_bit_math_h_l524_c3_4ef5_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node46_MUX_bit_math_h_l524_c3_4ef5_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node46_MUX_bit_math_h_l524_c3_4ef5_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node46_MUX_bit_math_h_l524_c3_4ef5_cond : unsigned(0 downto 0);
 variable VAR_layer0_node47 : unsigned(7 downto 0);
 variable VAR_layer0_node47_MUX_bit_math_h_l535_c3_21f3_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node47_MUX_bit_math_h_l535_c3_21f3_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node47_MUX_bit_math_h_l535_c3_21f3_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node47_MUX_bit_math_h_l535_c3_21f3_cond : unsigned(0 downto 0);
 variable VAR_layer0_node48 : unsigned(7 downto 0);
 variable VAR_layer0_node48_MUX_bit_math_h_l546_c3_5be4_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node48_MUX_bit_math_h_l546_c3_5be4_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node48_MUX_bit_math_h_l546_c3_5be4_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node48_MUX_bit_math_h_l546_c3_5be4_cond : unsigned(0 downto 0);
 variable VAR_layer0_node49 : unsigned(7 downto 0);
 variable VAR_layer0_node49_MUX_bit_math_h_l557_c3_3410_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node49_MUX_bit_math_h_l557_c3_3410_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node49_MUX_bit_math_h_l557_c3_3410_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node49_MUX_bit_math_h_l557_c3_3410_cond : unsigned(0 downto 0);
 variable VAR_layer0_node50 : unsigned(7 downto 0);
 variable VAR_layer0_node50_MUX_bit_math_h_l568_c3_4522_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node50_MUX_bit_math_h_l568_c3_4522_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node50_MUX_bit_math_h_l568_c3_4522_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node50_MUX_bit_math_h_l568_c3_4522_cond : unsigned(0 downto 0);
 variable VAR_layer0_node51 : unsigned(7 downto 0);
 variable VAR_layer0_node51_MUX_bit_math_h_l579_c3_8398_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node51_MUX_bit_math_h_l579_c3_8398_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node51_MUX_bit_math_h_l579_c3_8398_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node51_MUX_bit_math_h_l579_c3_8398_cond : unsigned(0 downto 0);
 variable VAR_layer0_node52 : unsigned(7 downto 0);
 variable VAR_layer0_node52_MUX_bit_math_h_l590_c3_6d3d_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node52_MUX_bit_math_h_l590_c3_6d3d_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node52_MUX_bit_math_h_l590_c3_6d3d_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node52_MUX_bit_math_h_l590_c3_6d3d_cond : unsigned(0 downto 0);
 variable VAR_layer0_node53 : unsigned(7 downto 0);
 variable VAR_layer0_node53_MUX_bit_math_h_l601_c3_6dc2_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node53_MUX_bit_math_h_l601_c3_6dc2_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node53_MUX_bit_math_h_l601_c3_6dc2_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node53_MUX_bit_math_h_l601_c3_6dc2_cond : unsigned(0 downto 0);
 variable VAR_layer0_node54 : unsigned(7 downto 0);
 variable VAR_layer0_node54_MUX_bit_math_h_l612_c3_cab9_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node54_MUX_bit_math_h_l612_c3_cab9_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node54_MUX_bit_math_h_l612_c3_cab9_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node54_MUX_bit_math_h_l612_c3_cab9_cond : unsigned(0 downto 0);
 variable VAR_layer0_node55 : unsigned(7 downto 0);
 variable VAR_layer0_node55_MUX_bit_math_h_l623_c3_2e5e_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node55_MUX_bit_math_h_l623_c3_2e5e_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node55_MUX_bit_math_h_l623_c3_2e5e_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node55_MUX_bit_math_h_l623_c3_2e5e_cond : unsigned(0 downto 0);
 variable VAR_layer0_node56 : unsigned(7 downto 0);
 variable VAR_layer0_node56_MUX_bit_math_h_l634_c3_ab19_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node56_MUX_bit_math_h_l634_c3_ab19_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node56_MUX_bit_math_h_l634_c3_ab19_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node56_MUX_bit_math_h_l634_c3_ab19_cond : unsigned(0 downto 0);
 variable VAR_layer0_node57 : unsigned(7 downto 0);
 variable VAR_layer0_node57_MUX_bit_math_h_l645_c3_cec5_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node57_MUX_bit_math_h_l645_c3_cec5_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node57_MUX_bit_math_h_l645_c3_cec5_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node57_MUX_bit_math_h_l645_c3_cec5_cond : unsigned(0 downto 0);
 variable VAR_layer0_node58 : unsigned(7 downto 0);
 variable VAR_layer0_node58_MUX_bit_math_h_l656_c3_312b_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node58_MUX_bit_math_h_l656_c3_312b_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node58_MUX_bit_math_h_l656_c3_312b_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node58_MUX_bit_math_h_l656_c3_312b_cond : unsigned(0 downto 0);
 variable VAR_layer0_node59 : unsigned(7 downto 0);
 variable VAR_layer0_node59_MUX_bit_math_h_l667_c3_672d_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node59_MUX_bit_math_h_l667_c3_672d_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node59_MUX_bit_math_h_l667_c3_672d_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node59_MUX_bit_math_h_l667_c3_672d_cond : unsigned(0 downto 0);
 variable VAR_layer0_node60 : unsigned(7 downto 0);
 variable VAR_layer0_node60_MUX_bit_math_h_l678_c3_9a42_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node60_MUX_bit_math_h_l678_c3_9a42_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node60_MUX_bit_math_h_l678_c3_9a42_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node60_MUX_bit_math_h_l678_c3_9a42_cond : unsigned(0 downto 0);
 variable VAR_layer0_node61 : unsigned(7 downto 0);
 variable VAR_layer0_node61_MUX_bit_math_h_l689_c3_be95_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node61_MUX_bit_math_h_l689_c3_be95_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node61_MUX_bit_math_h_l689_c3_be95_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node61_MUX_bit_math_h_l689_c3_be95_cond : unsigned(0 downto 0);
 variable VAR_layer0_node62 : unsigned(7 downto 0);
 variable VAR_layer0_node62_MUX_bit_math_h_l700_c3_8a98_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node62_MUX_bit_math_h_l700_c3_8a98_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node62_MUX_bit_math_h_l700_c3_8a98_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node62_MUX_bit_math_h_l700_c3_8a98_cond : unsigned(0 downto 0);
 variable VAR_layer0_node63 : unsigned(7 downto 0);
 variable VAR_layer0_node63_MUX_bit_math_h_l711_c3_45fc_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node63_MUX_bit_math_h_l711_c3_45fc_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node63_MUX_bit_math_h_l711_c3_45fc_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node63_MUX_bit_math_h_l711_c3_45fc_cond : unsigned(0 downto 0);
 variable VAR_sel1 : unsigned(0 downto 0);
 variable VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output : unsigned(0 downto 0);
 variable VAR_layer1_node0 : unsigned(7 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l728_c3_2ff0_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l728_c3_2ff0_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l728_c3_2ff0_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l728_c3_2ff0_cond : unsigned(0 downto 0);
 variable VAR_layer1_node1 : unsigned(7 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l739_c3_8d8d_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l739_c3_8d8d_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l739_c3_8d8d_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l739_c3_8d8d_cond : unsigned(0 downto 0);
 variable VAR_layer1_node2 : unsigned(7 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l750_c3_7ed6_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l750_c3_7ed6_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l750_c3_7ed6_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l750_c3_7ed6_cond : unsigned(0 downto 0);
 variable VAR_layer1_node3 : unsigned(7 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l761_c3_68af_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l761_c3_68af_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l761_c3_68af_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l761_c3_68af_cond : unsigned(0 downto 0);
 variable VAR_layer1_node4 : unsigned(7 downto 0);
 variable VAR_layer1_node4_MUX_bit_math_h_l772_c3_e8c5_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node4_MUX_bit_math_h_l772_c3_e8c5_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node4_MUX_bit_math_h_l772_c3_e8c5_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node4_MUX_bit_math_h_l772_c3_e8c5_cond : unsigned(0 downto 0);
 variable VAR_layer1_node5 : unsigned(7 downto 0);
 variable VAR_layer1_node5_MUX_bit_math_h_l783_c3_7ab9_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node5_MUX_bit_math_h_l783_c3_7ab9_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node5_MUX_bit_math_h_l783_c3_7ab9_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node5_MUX_bit_math_h_l783_c3_7ab9_cond : unsigned(0 downto 0);
 variable VAR_layer1_node6 : unsigned(7 downto 0);
 variable VAR_layer1_node6_MUX_bit_math_h_l794_c3_1dbe_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node6_MUX_bit_math_h_l794_c3_1dbe_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node6_MUX_bit_math_h_l794_c3_1dbe_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node6_MUX_bit_math_h_l794_c3_1dbe_cond : unsigned(0 downto 0);
 variable VAR_layer1_node7 : unsigned(7 downto 0);
 variable VAR_layer1_node7_MUX_bit_math_h_l805_c3_6dfe_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node7_MUX_bit_math_h_l805_c3_6dfe_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node7_MUX_bit_math_h_l805_c3_6dfe_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node7_MUX_bit_math_h_l805_c3_6dfe_cond : unsigned(0 downto 0);
 variable VAR_layer1_node8 : unsigned(7 downto 0);
 variable VAR_layer1_node8_MUX_bit_math_h_l816_c3_5d19_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node8_MUX_bit_math_h_l816_c3_5d19_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node8_MUX_bit_math_h_l816_c3_5d19_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node8_MUX_bit_math_h_l816_c3_5d19_cond : unsigned(0 downto 0);
 variable VAR_layer1_node9 : unsigned(7 downto 0);
 variable VAR_layer1_node9_MUX_bit_math_h_l827_c3_fe3d_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node9_MUX_bit_math_h_l827_c3_fe3d_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node9_MUX_bit_math_h_l827_c3_fe3d_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node9_MUX_bit_math_h_l827_c3_fe3d_cond : unsigned(0 downto 0);
 variable VAR_layer1_node10 : unsigned(7 downto 0);
 variable VAR_layer1_node10_MUX_bit_math_h_l838_c3_cc59_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node10_MUX_bit_math_h_l838_c3_cc59_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node10_MUX_bit_math_h_l838_c3_cc59_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node10_MUX_bit_math_h_l838_c3_cc59_cond : unsigned(0 downto 0);
 variable VAR_layer1_node11 : unsigned(7 downto 0);
 variable VAR_layer1_node11_MUX_bit_math_h_l849_c3_6ba8_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node11_MUX_bit_math_h_l849_c3_6ba8_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node11_MUX_bit_math_h_l849_c3_6ba8_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node11_MUX_bit_math_h_l849_c3_6ba8_cond : unsigned(0 downto 0);
 variable VAR_layer1_node12 : unsigned(7 downto 0);
 variable VAR_layer1_node12_MUX_bit_math_h_l860_c3_e057_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node12_MUX_bit_math_h_l860_c3_e057_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node12_MUX_bit_math_h_l860_c3_e057_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node12_MUX_bit_math_h_l860_c3_e057_cond : unsigned(0 downto 0);
 variable VAR_layer1_node13 : unsigned(7 downto 0);
 variable VAR_layer1_node13_MUX_bit_math_h_l871_c3_aad3_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node13_MUX_bit_math_h_l871_c3_aad3_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node13_MUX_bit_math_h_l871_c3_aad3_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node13_MUX_bit_math_h_l871_c3_aad3_cond : unsigned(0 downto 0);
 variable VAR_layer1_node14 : unsigned(7 downto 0);
 variable VAR_layer1_node14_MUX_bit_math_h_l882_c3_0d3c_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node14_MUX_bit_math_h_l882_c3_0d3c_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node14_MUX_bit_math_h_l882_c3_0d3c_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node14_MUX_bit_math_h_l882_c3_0d3c_cond : unsigned(0 downto 0);
 variable VAR_layer1_node15 : unsigned(7 downto 0);
 variable VAR_layer1_node15_MUX_bit_math_h_l893_c3_6301_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node15_MUX_bit_math_h_l893_c3_6301_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node15_MUX_bit_math_h_l893_c3_6301_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node15_MUX_bit_math_h_l893_c3_6301_cond : unsigned(0 downto 0);
 variable VAR_layer1_node16 : unsigned(7 downto 0);
 variable VAR_layer1_node16_MUX_bit_math_h_l904_c3_60f0_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node16_MUX_bit_math_h_l904_c3_60f0_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node16_MUX_bit_math_h_l904_c3_60f0_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node16_MUX_bit_math_h_l904_c3_60f0_cond : unsigned(0 downto 0);
 variable VAR_layer1_node17 : unsigned(7 downto 0);
 variable VAR_layer1_node17_MUX_bit_math_h_l915_c3_d47f_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node17_MUX_bit_math_h_l915_c3_d47f_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node17_MUX_bit_math_h_l915_c3_d47f_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node17_MUX_bit_math_h_l915_c3_d47f_cond : unsigned(0 downto 0);
 variable VAR_layer1_node18 : unsigned(7 downto 0);
 variable VAR_layer1_node18_MUX_bit_math_h_l926_c3_678f_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node18_MUX_bit_math_h_l926_c3_678f_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node18_MUX_bit_math_h_l926_c3_678f_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node18_MUX_bit_math_h_l926_c3_678f_cond : unsigned(0 downto 0);
 variable VAR_layer1_node19 : unsigned(7 downto 0);
 variable VAR_layer1_node19_MUX_bit_math_h_l937_c3_eb8f_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node19_MUX_bit_math_h_l937_c3_eb8f_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node19_MUX_bit_math_h_l937_c3_eb8f_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node19_MUX_bit_math_h_l937_c3_eb8f_cond : unsigned(0 downto 0);
 variable VAR_layer1_node20 : unsigned(7 downto 0);
 variable VAR_layer1_node20_MUX_bit_math_h_l948_c3_588a_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node20_MUX_bit_math_h_l948_c3_588a_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node20_MUX_bit_math_h_l948_c3_588a_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node20_MUX_bit_math_h_l948_c3_588a_cond : unsigned(0 downto 0);
 variable VAR_layer1_node21 : unsigned(7 downto 0);
 variable VAR_layer1_node21_MUX_bit_math_h_l959_c3_1823_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node21_MUX_bit_math_h_l959_c3_1823_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node21_MUX_bit_math_h_l959_c3_1823_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node21_MUX_bit_math_h_l959_c3_1823_cond : unsigned(0 downto 0);
 variable VAR_layer1_node22 : unsigned(7 downto 0);
 variable VAR_layer1_node22_MUX_bit_math_h_l970_c3_6904_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node22_MUX_bit_math_h_l970_c3_6904_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node22_MUX_bit_math_h_l970_c3_6904_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node22_MUX_bit_math_h_l970_c3_6904_cond : unsigned(0 downto 0);
 variable VAR_layer1_node23 : unsigned(7 downto 0);
 variable VAR_layer1_node23_MUX_bit_math_h_l981_c3_f890_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node23_MUX_bit_math_h_l981_c3_f890_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node23_MUX_bit_math_h_l981_c3_f890_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node23_MUX_bit_math_h_l981_c3_f890_cond : unsigned(0 downto 0);
 variable VAR_layer1_node24 : unsigned(7 downto 0);
 variable VAR_layer1_node24_MUX_bit_math_h_l992_c3_4e65_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node24_MUX_bit_math_h_l992_c3_4e65_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node24_MUX_bit_math_h_l992_c3_4e65_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node24_MUX_bit_math_h_l992_c3_4e65_cond : unsigned(0 downto 0);
 variable VAR_layer1_node25 : unsigned(7 downto 0);
 variable VAR_layer1_node25_MUX_bit_math_h_l1003_c3_f943_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node25_MUX_bit_math_h_l1003_c3_f943_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node25_MUX_bit_math_h_l1003_c3_f943_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node25_MUX_bit_math_h_l1003_c3_f943_cond : unsigned(0 downto 0);
 variable VAR_layer1_node26 : unsigned(7 downto 0);
 variable VAR_layer1_node26_MUX_bit_math_h_l1014_c3_aa20_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node26_MUX_bit_math_h_l1014_c3_aa20_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node26_MUX_bit_math_h_l1014_c3_aa20_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node26_MUX_bit_math_h_l1014_c3_aa20_cond : unsigned(0 downto 0);
 variable VAR_layer1_node27 : unsigned(7 downto 0);
 variable VAR_layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_cond : unsigned(0 downto 0);
 variable VAR_layer1_node28 : unsigned(7 downto 0);
 variable VAR_layer1_node28_MUX_bit_math_h_l1036_c3_85a0_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node28_MUX_bit_math_h_l1036_c3_85a0_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node28_MUX_bit_math_h_l1036_c3_85a0_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node28_MUX_bit_math_h_l1036_c3_85a0_cond : unsigned(0 downto 0);
 variable VAR_layer1_node29 : unsigned(7 downto 0);
 variable VAR_layer1_node29_MUX_bit_math_h_l1047_c3_953f_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node29_MUX_bit_math_h_l1047_c3_953f_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node29_MUX_bit_math_h_l1047_c3_953f_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node29_MUX_bit_math_h_l1047_c3_953f_cond : unsigned(0 downto 0);
 variable VAR_layer1_node30 : unsigned(7 downto 0);
 variable VAR_layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_cond : unsigned(0 downto 0);
 variable VAR_layer1_node31 : unsigned(7 downto 0);
 variable VAR_layer1_node31_MUX_bit_math_h_l1069_c3_82fc_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node31_MUX_bit_math_h_l1069_c3_82fc_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node31_MUX_bit_math_h_l1069_c3_82fc_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node31_MUX_bit_math_h_l1069_c3_82fc_cond : unsigned(0 downto 0);
 variable VAR_sel2 : unsigned(0 downto 0);
 variable VAR_uint7_2_2_bit_math_h_l1082_c10_12df_return_output : unsigned(0 downto 0);
 variable VAR_layer2_node0 : unsigned(7 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l1086_c3_4e60_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l1086_c3_4e60_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l1086_c3_4e60_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l1086_c3_4e60_cond : unsigned(0 downto 0);
 variable VAR_layer2_node1 : unsigned(7 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l1097_c3_12bb_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l1097_c3_12bb_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l1097_c3_12bb_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l1097_c3_12bb_cond : unsigned(0 downto 0);
 variable VAR_layer2_node2 : unsigned(7 downto 0);
 variable VAR_layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_cond : unsigned(0 downto 0);
 variable VAR_layer2_node3 : unsigned(7 downto 0);
 variable VAR_layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_cond : unsigned(0 downto 0);
 variable VAR_layer2_node4 : unsigned(7 downto 0);
 variable VAR_layer2_node4_MUX_bit_math_h_l1130_c3_3de0_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node4_MUX_bit_math_h_l1130_c3_3de0_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node4_MUX_bit_math_h_l1130_c3_3de0_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node4_MUX_bit_math_h_l1130_c3_3de0_cond : unsigned(0 downto 0);
 variable VAR_layer2_node5 : unsigned(7 downto 0);
 variable VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_cond : unsigned(0 downto 0);
 variable VAR_layer2_node6 : unsigned(7 downto 0);
 variable VAR_layer2_node6_MUX_bit_math_h_l1152_c3_3828_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node6_MUX_bit_math_h_l1152_c3_3828_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node6_MUX_bit_math_h_l1152_c3_3828_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node6_MUX_bit_math_h_l1152_c3_3828_cond : unsigned(0 downto 0);
 variable VAR_layer2_node7 : unsigned(7 downto 0);
 variable VAR_layer2_node7_MUX_bit_math_h_l1163_c3_f226_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node7_MUX_bit_math_h_l1163_c3_f226_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node7_MUX_bit_math_h_l1163_c3_f226_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node7_MUX_bit_math_h_l1163_c3_f226_cond : unsigned(0 downto 0);
 variable VAR_layer2_node8 : unsigned(7 downto 0);
 variable VAR_layer2_node8_MUX_bit_math_h_l1174_c3_49b7_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node8_MUX_bit_math_h_l1174_c3_49b7_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node8_MUX_bit_math_h_l1174_c3_49b7_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node8_MUX_bit_math_h_l1174_c3_49b7_cond : unsigned(0 downto 0);
 variable VAR_layer2_node9 : unsigned(7 downto 0);
 variable VAR_layer2_node9_MUX_bit_math_h_l1185_c3_934f_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node9_MUX_bit_math_h_l1185_c3_934f_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node9_MUX_bit_math_h_l1185_c3_934f_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node9_MUX_bit_math_h_l1185_c3_934f_cond : unsigned(0 downto 0);
 variable VAR_layer2_node10 : unsigned(7 downto 0);
 variable VAR_layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_cond : unsigned(0 downto 0);
 variable VAR_layer2_node11 : unsigned(7 downto 0);
 variable VAR_layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_cond : unsigned(0 downto 0);
 variable VAR_layer2_node12 : unsigned(7 downto 0);
 variable VAR_layer2_node12_MUX_bit_math_h_l1218_c3_0726_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node12_MUX_bit_math_h_l1218_c3_0726_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node12_MUX_bit_math_h_l1218_c3_0726_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node12_MUX_bit_math_h_l1218_c3_0726_cond : unsigned(0 downto 0);
 variable VAR_layer2_node13 : unsigned(7 downto 0);
 variable VAR_layer2_node13_MUX_bit_math_h_l1229_c3_754d_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node13_MUX_bit_math_h_l1229_c3_754d_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node13_MUX_bit_math_h_l1229_c3_754d_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node13_MUX_bit_math_h_l1229_c3_754d_cond : unsigned(0 downto 0);
 variable VAR_layer2_node14 : unsigned(7 downto 0);
 variable VAR_layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_cond : unsigned(0 downto 0);
 variable VAR_layer2_node15 : unsigned(7 downto 0);
 variable VAR_layer2_node15_MUX_bit_math_h_l1251_c3_57b2_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node15_MUX_bit_math_h_l1251_c3_57b2_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node15_MUX_bit_math_h_l1251_c3_57b2_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node15_MUX_bit_math_h_l1251_c3_57b2_cond : unsigned(0 downto 0);
 variable VAR_sel3 : unsigned(0 downto 0);
 variable VAR_uint7_3_3_bit_math_h_l1264_c10_4cf0_return_output : unsigned(0 downto 0);
 variable VAR_layer3_node0 : unsigned(7 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_cond : unsigned(0 downto 0);
 variable VAR_layer3_node1 : unsigned(7 downto 0);
 variable VAR_layer3_node1_MUX_bit_math_h_l1279_c3_73ae_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node1_MUX_bit_math_h_l1279_c3_73ae_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node1_MUX_bit_math_h_l1279_c3_73ae_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node1_MUX_bit_math_h_l1279_c3_73ae_cond : unsigned(0 downto 0);
 variable VAR_layer3_node2 : unsigned(7 downto 0);
 variable VAR_layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_cond : unsigned(0 downto 0);
 variable VAR_layer3_node3 : unsigned(7 downto 0);
 variable VAR_layer3_node3_MUX_bit_math_h_l1301_c3_827d_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node3_MUX_bit_math_h_l1301_c3_827d_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node3_MUX_bit_math_h_l1301_c3_827d_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node3_MUX_bit_math_h_l1301_c3_827d_cond : unsigned(0 downto 0);
 variable VAR_layer3_node4 : unsigned(7 downto 0);
 variable VAR_layer3_node4_MUX_bit_math_h_l1312_c3_ca04_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node4_MUX_bit_math_h_l1312_c3_ca04_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node4_MUX_bit_math_h_l1312_c3_ca04_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node4_MUX_bit_math_h_l1312_c3_ca04_cond : unsigned(0 downto 0);
 variable VAR_layer3_node5 : unsigned(7 downto 0);
 variable VAR_layer3_node5_MUX_bit_math_h_l1323_c3_56dd_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node5_MUX_bit_math_h_l1323_c3_56dd_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node5_MUX_bit_math_h_l1323_c3_56dd_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node5_MUX_bit_math_h_l1323_c3_56dd_cond : unsigned(0 downto 0);
 variable VAR_layer3_node6 : unsigned(7 downto 0);
 variable VAR_layer3_node6_MUX_bit_math_h_l1334_c3_07bd_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node6_MUX_bit_math_h_l1334_c3_07bd_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node6_MUX_bit_math_h_l1334_c3_07bd_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node6_MUX_bit_math_h_l1334_c3_07bd_cond : unsigned(0 downto 0);
 variable VAR_layer3_node7 : unsigned(7 downto 0);
 variable VAR_layer3_node7_MUX_bit_math_h_l1345_c3_5a50_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node7_MUX_bit_math_h_l1345_c3_5a50_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node7_MUX_bit_math_h_l1345_c3_5a50_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node7_MUX_bit_math_h_l1345_c3_5a50_cond : unsigned(0 downto 0);
 variable VAR_sel4 : unsigned(0 downto 0);
 variable VAR_uint7_4_4_bit_math_h_l1358_c10_0af5_return_output : unsigned(0 downto 0);
 variable VAR_layer4_node0 : unsigned(7 downto 0);
 variable VAR_layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_iftrue : unsigned(7 downto 0);
 variable VAR_layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_iffalse : unsigned(7 downto 0);
 variable VAR_layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_return_output : unsigned(7 downto 0);
 variable VAR_layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_cond : unsigned(0 downto 0);
 variable VAR_layer4_node1 : unsigned(7 downto 0);
 variable VAR_layer4_node1_MUX_bit_math_h_l1373_c3_402b_iftrue : unsigned(7 downto 0);
 variable VAR_layer4_node1_MUX_bit_math_h_l1373_c3_402b_iffalse : unsigned(7 downto 0);
 variable VAR_layer4_node1_MUX_bit_math_h_l1373_c3_402b_return_output : unsigned(7 downto 0);
 variable VAR_layer4_node1_MUX_bit_math_h_l1373_c3_402b_cond : unsigned(0 downto 0);
 variable VAR_layer4_node2 : unsigned(7 downto 0);
 variable VAR_layer4_node2_MUX_bit_math_h_l1384_c3_5f80_iftrue : unsigned(7 downto 0);
 variable VAR_layer4_node2_MUX_bit_math_h_l1384_c3_5f80_iffalse : unsigned(7 downto 0);
 variable VAR_layer4_node2_MUX_bit_math_h_l1384_c3_5f80_return_output : unsigned(7 downto 0);
 variable VAR_layer4_node2_MUX_bit_math_h_l1384_c3_5f80_cond : unsigned(0 downto 0);
 variable VAR_layer4_node3 : unsigned(7 downto 0);
 variable VAR_layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_iftrue : unsigned(7 downto 0);
 variable VAR_layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_iffalse : unsigned(7 downto 0);
 variable VAR_layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_return_output : unsigned(7 downto 0);
 variable VAR_layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_cond : unsigned(0 downto 0);
 variable VAR_sel5 : unsigned(0 downto 0);
 variable VAR_uint7_5_5_bit_math_h_l1408_c10_41c5_return_output : unsigned(0 downto 0);
 variable VAR_layer5_node0 : unsigned(7 downto 0);
 variable VAR_layer5_node0_MUX_bit_math_h_l1412_c3_19e3_iftrue : unsigned(7 downto 0);
 variable VAR_layer5_node0_MUX_bit_math_h_l1412_c3_19e3_iffalse : unsigned(7 downto 0);
 variable VAR_layer5_node0_MUX_bit_math_h_l1412_c3_19e3_return_output : unsigned(7 downto 0);
 variable VAR_layer5_node0_MUX_bit_math_h_l1412_c3_19e3_cond : unsigned(0 downto 0);
 variable VAR_layer5_node1 : unsigned(7 downto 0);
 variable VAR_layer5_node1_MUX_bit_math_h_l1423_c3_11f1_iftrue : unsigned(7 downto 0);
 variable VAR_layer5_node1_MUX_bit_math_h_l1423_c3_11f1_iffalse : unsigned(7 downto 0);
 variable VAR_layer5_node1_MUX_bit_math_h_l1423_c3_11f1_return_output : unsigned(7 downto 0);
 variable VAR_layer5_node1_MUX_bit_math_h_l1423_c3_11f1_cond : unsigned(0 downto 0);
 variable VAR_sel6 : unsigned(0 downto 0);
 variable VAR_uint7_6_6_bit_math_h_l1436_c10_c6df_return_output : unsigned(0 downto 0);
 variable VAR_layer6_node0 : unsigned(7 downto 0);
 variable VAR_layer6_node0_MUX_bit_math_h_l1440_c3_f906_iftrue : unsigned(7 downto 0);
 variable VAR_layer6_node0_MUX_bit_math_h_l1440_c3_f906_iffalse : unsigned(7 downto 0);
 variable VAR_layer6_node0_MUX_bit_math_h_l1440_c3_f906_return_output : unsigned(7 downto 0);
 variable VAR_layer6_node0_MUX_bit_math_h_l1440_c3_f906_cond : unsigned(0 downto 0);
begin

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_sel := sel;
     VAR_in0 := in0;
     VAR_in1 := in1;
     VAR_in2 := in2;
     VAR_in3 := in3;
     VAR_in4 := in4;
     VAR_in5 := in5;
     VAR_in6 := in6;
     VAR_in7 := in7;
     VAR_in8 := in8;
     VAR_in9 := in9;
     VAR_in10 := in10;
     VAR_in11 := in11;
     VAR_in12 := in12;
     VAR_in13 := in13;
     VAR_in14 := in14;
     VAR_in15 := in15;
     VAR_in16 := in16;
     VAR_in17 := in17;
     VAR_in18 := in18;
     VAR_in19 := in19;
     VAR_in20 := in20;
     VAR_in21 := in21;
     VAR_in22 := in22;
     VAR_in23 := in23;
     VAR_in24 := in24;
     VAR_in25 := in25;
     VAR_in26 := in26;
     VAR_in27 := in27;
     VAR_in28 := in28;
     VAR_in29 := in29;
     VAR_in30 := in30;
     VAR_in31 := in31;
     VAR_in32 := in32;
     VAR_in33 := in33;
     VAR_in34 := in34;
     VAR_in35 := in35;
     VAR_in36 := in36;
     VAR_in37 := in37;
     VAR_in38 := in38;
     VAR_in39 := in39;
     VAR_in40 := in40;
     VAR_in41 := in41;
     VAR_in42 := in42;
     VAR_in43 := in43;
     VAR_in44 := in44;
     VAR_in45 := in45;
     VAR_in46 := in46;
     VAR_in47 := in47;
     VAR_in48 := in48;
     VAR_in49 := in49;
     VAR_in50 := in50;
     VAR_in51 := in51;
     VAR_in52 := in52;
     VAR_in53 := in53;
     VAR_in54 := in54;
     VAR_in55 := in55;
     VAR_in56 := in56;
     VAR_in57 := in57;
     VAR_in58 := in58;
     VAR_in59 := in59;
     VAR_in60 := in60;
     VAR_in61 := in61;
     VAR_in62 := in62;
     VAR_in63 := in63;
     VAR_in64 := in64;
     VAR_in65 := in65;
     VAR_in66 := in66;
     VAR_in67 := in67;
     VAR_in68 := in68;
     VAR_in69 := in69;
     VAR_in70 := in70;
     VAR_in71 := in71;
     VAR_in72 := in72;
     VAR_in73 := in73;
     VAR_in74 := in74;
     VAR_in75 := in75;
     VAR_in76 := in76;
     VAR_in77 := in77;
     VAR_in78 := in78;
     VAR_in79 := in79;
     VAR_in80 := in80;
     VAR_in81 := in81;
     VAR_in82 := in82;
     VAR_in83 := in83;
     VAR_in84 := in84;
     VAR_in85 := in85;
     VAR_in86 := in86;
     VAR_in87 := in87;
     VAR_in88 := in88;
     VAR_in89 := in89;
     VAR_in90 := in90;
     VAR_in91 := in91;
     VAR_in92 := in92;
     VAR_in93 := in93;
     VAR_in94 := in94;
     VAR_in95 := in95;
     VAR_in96 := in96;
     VAR_in97 := in97;
     VAR_in98 := in98;
     VAR_in99 := in99;
     VAR_in100 := in100;
     VAR_in101 := in101;
     VAR_in102 := in102;
     VAR_in103 := in103;
     VAR_in104 := in104;
     VAR_in105 := in105;
     VAR_in106 := in106;
     VAR_in107 := in107;
     VAR_in108 := in108;
     VAR_in109 := in109;
     VAR_in110 := in110;
     VAR_in111 := in111;
     VAR_in112 := in112;
     VAR_in113 := in113;
     VAR_in114 := in114;
     VAR_in115 := in115;
     VAR_in116 := in116;
     VAR_in117 := in117;
     VAR_in118 := in118;
     VAR_in119 := in119;
     VAR_in120 := in120;
     VAR_in121 := in121;
     VAR_in122 := in122;
     VAR_in123 := in123;
     VAR_in124 := in124;
     VAR_in125 := in125;
     VAR_in126 := in126;
     VAR_in127 := in127;

     -- Submodule level 0
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_5c06_iffalse := VAR_in0;
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_5c06_iftrue := VAR_in1;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_282b_iffalse := VAR_in10;
     VAR_layer0_node50_MUX_bit_math_h_l568_c3_4522_iffalse := VAR_in100;
     VAR_layer0_node50_MUX_bit_math_h_l568_c3_4522_iftrue := VAR_in101;
     VAR_layer0_node51_MUX_bit_math_h_l579_c3_8398_iffalse := VAR_in102;
     VAR_layer0_node51_MUX_bit_math_h_l579_c3_8398_iftrue := VAR_in103;
     VAR_layer0_node52_MUX_bit_math_h_l590_c3_6d3d_iffalse := VAR_in104;
     VAR_layer0_node52_MUX_bit_math_h_l590_c3_6d3d_iftrue := VAR_in105;
     VAR_layer0_node53_MUX_bit_math_h_l601_c3_6dc2_iffalse := VAR_in106;
     VAR_layer0_node53_MUX_bit_math_h_l601_c3_6dc2_iftrue := VAR_in107;
     VAR_layer0_node54_MUX_bit_math_h_l612_c3_cab9_iffalse := VAR_in108;
     VAR_layer0_node54_MUX_bit_math_h_l612_c3_cab9_iftrue := VAR_in109;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_282b_iftrue := VAR_in11;
     VAR_layer0_node55_MUX_bit_math_h_l623_c3_2e5e_iffalse := VAR_in110;
     VAR_layer0_node55_MUX_bit_math_h_l623_c3_2e5e_iftrue := VAR_in111;
     VAR_layer0_node56_MUX_bit_math_h_l634_c3_ab19_iffalse := VAR_in112;
     VAR_layer0_node56_MUX_bit_math_h_l634_c3_ab19_iftrue := VAR_in113;
     VAR_layer0_node57_MUX_bit_math_h_l645_c3_cec5_iffalse := VAR_in114;
     VAR_layer0_node57_MUX_bit_math_h_l645_c3_cec5_iftrue := VAR_in115;
     VAR_layer0_node58_MUX_bit_math_h_l656_c3_312b_iffalse := VAR_in116;
     VAR_layer0_node58_MUX_bit_math_h_l656_c3_312b_iftrue := VAR_in117;
     VAR_layer0_node59_MUX_bit_math_h_l667_c3_672d_iffalse := VAR_in118;
     VAR_layer0_node59_MUX_bit_math_h_l667_c3_672d_iftrue := VAR_in119;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_62f1_iffalse := VAR_in12;
     VAR_layer0_node60_MUX_bit_math_h_l678_c3_9a42_iffalse := VAR_in120;
     VAR_layer0_node60_MUX_bit_math_h_l678_c3_9a42_iftrue := VAR_in121;
     VAR_layer0_node61_MUX_bit_math_h_l689_c3_be95_iffalse := VAR_in122;
     VAR_layer0_node61_MUX_bit_math_h_l689_c3_be95_iftrue := VAR_in123;
     VAR_layer0_node62_MUX_bit_math_h_l700_c3_8a98_iffalse := VAR_in124;
     VAR_layer0_node62_MUX_bit_math_h_l700_c3_8a98_iftrue := VAR_in125;
     VAR_layer0_node63_MUX_bit_math_h_l711_c3_45fc_iffalse := VAR_in126;
     VAR_layer0_node63_MUX_bit_math_h_l711_c3_45fc_iftrue := VAR_in127;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_62f1_iftrue := VAR_in13;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_567b_iffalse := VAR_in14;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_567b_iftrue := VAR_in15;
     VAR_layer0_node8_MUX_bit_math_h_l106_c3_47e5_iffalse := VAR_in16;
     VAR_layer0_node8_MUX_bit_math_h_l106_c3_47e5_iftrue := VAR_in17;
     VAR_layer0_node9_MUX_bit_math_h_l117_c3_f097_iffalse := VAR_in18;
     VAR_layer0_node9_MUX_bit_math_h_l117_c3_f097_iftrue := VAR_in19;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_fa46_iffalse := VAR_in2;
     VAR_layer0_node10_MUX_bit_math_h_l128_c3_0e6c_iffalse := VAR_in20;
     VAR_layer0_node10_MUX_bit_math_h_l128_c3_0e6c_iftrue := VAR_in21;
     VAR_layer0_node11_MUX_bit_math_h_l139_c3_3ab9_iffalse := VAR_in22;
     VAR_layer0_node11_MUX_bit_math_h_l139_c3_3ab9_iftrue := VAR_in23;
     VAR_layer0_node12_MUX_bit_math_h_l150_c3_e611_iffalse := VAR_in24;
     VAR_layer0_node12_MUX_bit_math_h_l150_c3_e611_iftrue := VAR_in25;
     VAR_layer0_node13_MUX_bit_math_h_l161_c3_e037_iffalse := VAR_in26;
     VAR_layer0_node13_MUX_bit_math_h_l161_c3_e037_iftrue := VAR_in27;
     VAR_layer0_node14_MUX_bit_math_h_l172_c3_ad25_iffalse := VAR_in28;
     VAR_layer0_node14_MUX_bit_math_h_l172_c3_ad25_iftrue := VAR_in29;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_fa46_iftrue := VAR_in3;
     VAR_layer0_node15_MUX_bit_math_h_l183_c3_dacd_iffalse := VAR_in30;
     VAR_layer0_node15_MUX_bit_math_h_l183_c3_dacd_iftrue := VAR_in31;
     VAR_layer0_node16_MUX_bit_math_h_l194_c3_5393_iffalse := VAR_in32;
     VAR_layer0_node16_MUX_bit_math_h_l194_c3_5393_iftrue := VAR_in33;
     VAR_layer0_node17_MUX_bit_math_h_l205_c3_4246_iffalse := VAR_in34;
     VAR_layer0_node17_MUX_bit_math_h_l205_c3_4246_iftrue := VAR_in35;
     VAR_layer0_node18_MUX_bit_math_h_l216_c3_2748_iffalse := VAR_in36;
     VAR_layer0_node18_MUX_bit_math_h_l216_c3_2748_iftrue := VAR_in37;
     VAR_layer0_node19_MUX_bit_math_h_l227_c3_1dae_iffalse := VAR_in38;
     VAR_layer0_node19_MUX_bit_math_h_l227_c3_1dae_iftrue := VAR_in39;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_f68a_iffalse := VAR_in4;
     VAR_layer0_node20_MUX_bit_math_h_l238_c3_e7c7_iffalse := VAR_in40;
     VAR_layer0_node20_MUX_bit_math_h_l238_c3_e7c7_iftrue := VAR_in41;
     VAR_layer0_node21_MUX_bit_math_h_l249_c3_8f8c_iffalse := VAR_in42;
     VAR_layer0_node21_MUX_bit_math_h_l249_c3_8f8c_iftrue := VAR_in43;
     VAR_layer0_node22_MUX_bit_math_h_l260_c3_321e_iffalse := VAR_in44;
     VAR_layer0_node22_MUX_bit_math_h_l260_c3_321e_iftrue := VAR_in45;
     VAR_layer0_node23_MUX_bit_math_h_l271_c3_86c3_iffalse := VAR_in46;
     VAR_layer0_node23_MUX_bit_math_h_l271_c3_86c3_iftrue := VAR_in47;
     VAR_layer0_node24_MUX_bit_math_h_l282_c3_2992_iffalse := VAR_in48;
     VAR_layer0_node24_MUX_bit_math_h_l282_c3_2992_iftrue := VAR_in49;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_f68a_iftrue := VAR_in5;
     VAR_layer0_node25_MUX_bit_math_h_l293_c3_ece2_iffalse := VAR_in50;
     VAR_layer0_node25_MUX_bit_math_h_l293_c3_ece2_iftrue := VAR_in51;
     VAR_layer0_node26_MUX_bit_math_h_l304_c3_7f9b_iffalse := VAR_in52;
     VAR_layer0_node26_MUX_bit_math_h_l304_c3_7f9b_iftrue := VAR_in53;
     VAR_layer0_node27_MUX_bit_math_h_l315_c3_5c0f_iffalse := VAR_in54;
     VAR_layer0_node27_MUX_bit_math_h_l315_c3_5c0f_iftrue := VAR_in55;
     VAR_layer0_node28_MUX_bit_math_h_l326_c3_12a3_iffalse := VAR_in56;
     VAR_layer0_node28_MUX_bit_math_h_l326_c3_12a3_iftrue := VAR_in57;
     VAR_layer0_node29_MUX_bit_math_h_l337_c3_cbb8_iffalse := VAR_in58;
     VAR_layer0_node29_MUX_bit_math_h_l337_c3_cbb8_iftrue := VAR_in59;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_b336_iffalse := VAR_in6;
     VAR_layer0_node30_MUX_bit_math_h_l348_c3_8c5c_iffalse := VAR_in60;
     VAR_layer0_node30_MUX_bit_math_h_l348_c3_8c5c_iftrue := VAR_in61;
     VAR_layer0_node31_MUX_bit_math_h_l359_c3_d6b9_iffalse := VAR_in62;
     VAR_layer0_node31_MUX_bit_math_h_l359_c3_d6b9_iftrue := VAR_in63;
     VAR_layer0_node32_MUX_bit_math_h_l370_c3_3d24_iffalse := VAR_in64;
     VAR_layer0_node32_MUX_bit_math_h_l370_c3_3d24_iftrue := VAR_in65;
     VAR_layer0_node33_MUX_bit_math_h_l381_c3_bdd0_iffalse := VAR_in66;
     VAR_layer0_node33_MUX_bit_math_h_l381_c3_bdd0_iftrue := VAR_in67;
     VAR_layer0_node34_MUX_bit_math_h_l392_c3_f617_iffalse := VAR_in68;
     VAR_layer0_node34_MUX_bit_math_h_l392_c3_f617_iftrue := VAR_in69;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_b336_iftrue := VAR_in7;
     VAR_layer0_node35_MUX_bit_math_h_l403_c3_683e_iffalse := VAR_in70;
     VAR_layer0_node35_MUX_bit_math_h_l403_c3_683e_iftrue := VAR_in71;
     VAR_layer0_node36_MUX_bit_math_h_l414_c3_cd2c_iffalse := VAR_in72;
     VAR_layer0_node36_MUX_bit_math_h_l414_c3_cd2c_iftrue := VAR_in73;
     VAR_layer0_node37_MUX_bit_math_h_l425_c3_2485_iffalse := VAR_in74;
     VAR_layer0_node37_MUX_bit_math_h_l425_c3_2485_iftrue := VAR_in75;
     VAR_layer0_node38_MUX_bit_math_h_l436_c3_c940_iffalse := VAR_in76;
     VAR_layer0_node38_MUX_bit_math_h_l436_c3_c940_iftrue := VAR_in77;
     VAR_layer0_node39_MUX_bit_math_h_l447_c3_b150_iffalse := VAR_in78;
     VAR_layer0_node39_MUX_bit_math_h_l447_c3_b150_iftrue := VAR_in79;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_07e7_iffalse := VAR_in8;
     VAR_layer0_node40_MUX_bit_math_h_l458_c3_c977_iffalse := VAR_in80;
     VAR_layer0_node40_MUX_bit_math_h_l458_c3_c977_iftrue := VAR_in81;
     VAR_layer0_node41_MUX_bit_math_h_l469_c3_b3bf_iffalse := VAR_in82;
     VAR_layer0_node41_MUX_bit_math_h_l469_c3_b3bf_iftrue := VAR_in83;
     VAR_layer0_node42_MUX_bit_math_h_l480_c3_c677_iffalse := VAR_in84;
     VAR_layer0_node42_MUX_bit_math_h_l480_c3_c677_iftrue := VAR_in85;
     VAR_layer0_node43_MUX_bit_math_h_l491_c3_2838_iffalse := VAR_in86;
     VAR_layer0_node43_MUX_bit_math_h_l491_c3_2838_iftrue := VAR_in87;
     VAR_layer0_node44_MUX_bit_math_h_l502_c3_6b96_iffalse := VAR_in88;
     VAR_layer0_node44_MUX_bit_math_h_l502_c3_6b96_iftrue := VAR_in89;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_07e7_iftrue := VAR_in9;
     VAR_layer0_node45_MUX_bit_math_h_l513_c3_b86e_iffalse := VAR_in90;
     VAR_layer0_node45_MUX_bit_math_h_l513_c3_b86e_iftrue := VAR_in91;
     VAR_layer0_node46_MUX_bit_math_h_l524_c3_4ef5_iffalse := VAR_in92;
     VAR_layer0_node46_MUX_bit_math_h_l524_c3_4ef5_iftrue := VAR_in93;
     VAR_layer0_node47_MUX_bit_math_h_l535_c3_21f3_iffalse := VAR_in94;
     VAR_layer0_node47_MUX_bit_math_h_l535_c3_21f3_iftrue := VAR_in95;
     VAR_layer0_node48_MUX_bit_math_h_l546_c3_5be4_iffalse := VAR_in96;
     VAR_layer0_node48_MUX_bit_math_h_l546_c3_5be4_iftrue := VAR_in97;
     VAR_layer0_node49_MUX_bit_math_h_l557_c3_3410_iffalse := VAR_in98;
     VAR_layer0_node49_MUX_bit_math_h_l557_c3_3410_iftrue := VAR_in99;
     -- uint7_1_1[bit_math_h_l724_c10_7c0a] LATENCY=0
     VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output := uint7_1_1(
     VAR_sel);

     -- uint7_3_3[bit_math_h_l1264_c10_4cf0] LATENCY=0
     VAR_uint7_3_3_bit_math_h_l1264_c10_4cf0_return_output := uint7_3_3(
     VAR_sel);

     -- uint7_2_2[bit_math_h_l1082_c10_12df] LATENCY=0
     VAR_uint7_2_2_bit_math_h_l1082_c10_12df_return_output := uint7_2_2(
     VAR_sel);

     -- uint7_0_0[bit_math_h_l14_c10_592f] LATENCY=0
     VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output := uint7_0_0(
     VAR_sel);

     -- uint7_5_5[bit_math_h_l1408_c10_41c5] LATENCY=0
     VAR_uint7_5_5_bit_math_h_l1408_c10_41c5_return_output := uint7_5_5(
     VAR_sel);

     -- uint7_6_6[bit_math_h_l1436_c10_c6df] LATENCY=0
     VAR_uint7_6_6_bit_math_h_l1436_c10_c6df_return_output := uint7_6_6(
     VAR_sel);

     -- uint7_4_4[bit_math_h_l1358_c10_0af5] LATENCY=0
     VAR_uint7_4_4_bit_math_h_l1358_c10_0af5_return_output := uint7_4_4(
     VAR_sel);

     -- Submodule level 1
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_5c06_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node10_MUX_bit_math_h_l128_c3_0e6c_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node11_MUX_bit_math_h_l139_c3_3ab9_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node12_MUX_bit_math_h_l150_c3_e611_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node13_MUX_bit_math_h_l161_c3_e037_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node14_MUX_bit_math_h_l172_c3_ad25_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node15_MUX_bit_math_h_l183_c3_dacd_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node16_MUX_bit_math_h_l194_c3_5393_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node17_MUX_bit_math_h_l205_c3_4246_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node18_MUX_bit_math_h_l216_c3_2748_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node19_MUX_bit_math_h_l227_c3_1dae_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_fa46_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node20_MUX_bit_math_h_l238_c3_e7c7_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node21_MUX_bit_math_h_l249_c3_8f8c_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node22_MUX_bit_math_h_l260_c3_321e_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node23_MUX_bit_math_h_l271_c3_86c3_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node24_MUX_bit_math_h_l282_c3_2992_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node25_MUX_bit_math_h_l293_c3_ece2_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node26_MUX_bit_math_h_l304_c3_7f9b_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node27_MUX_bit_math_h_l315_c3_5c0f_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node28_MUX_bit_math_h_l326_c3_12a3_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node29_MUX_bit_math_h_l337_c3_cbb8_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_f68a_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node30_MUX_bit_math_h_l348_c3_8c5c_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node31_MUX_bit_math_h_l359_c3_d6b9_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node32_MUX_bit_math_h_l370_c3_3d24_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node33_MUX_bit_math_h_l381_c3_bdd0_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node34_MUX_bit_math_h_l392_c3_f617_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node35_MUX_bit_math_h_l403_c3_683e_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node36_MUX_bit_math_h_l414_c3_cd2c_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node37_MUX_bit_math_h_l425_c3_2485_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node38_MUX_bit_math_h_l436_c3_c940_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node39_MUX_bit_math_h_l447_c3_b150_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_b336_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node40_MUX_bit_math_h_l458_c3_c977_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node41_MUX_bit_math_h_l469_c3_b3bf_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node42_MUX_bit_math_h_l480_c3_c677_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node43_MUX_bit_math_h_l491_c3_2838_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node44_MUX_bit_math_h_l502_c3_6b96_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node45_MUX_bit_math_h_l513_c3_b86e_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node46_MUX_bit_math_h_l524_c3_4ef5_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node47_MUX_bit_math_h_l535_c3_21f3_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node48_MUX_bit_math_h_l546_c3_5be4_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node49_MUX_bit_math_h_l557_c3_3410_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_07e7_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node50_MUX_bit_math_h_l568_c3_4522_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node51_MUX_bit_math_h_l579_c3_8398_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node52_MUX_bit_math_h_l590_c3_6d3d_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node53_MUX_bit_math_h_l601_c3_6dc2_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node54_MUX_bit_math_h_l612_c3_cab9_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node55_MUX_bit_math_h_l623_c3_2e5e_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node56_MUX_bit_math_h_l634_c3_ab19_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node57_MUX_bit_math_h_l645_c3_cec5_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node58_MUX_bit_math_h_l656_c3_312b_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node59_MUX_bit_math_h_l667_c3_672d_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_282b_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node60_MUX_bit_math_h_l678_c3_9a42_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node61_MUX_bit_math_h_l689_c3_be95_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node62_MUX_bit_math_h_l700_c3_8a98_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node63_MUX_bit_math_h_l711_c3_45fc_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_62f1_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_567b_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node8_MUX_bit_math_h_l106_c3_47e5_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer0_node9_MUX_bit_math_h_l117_c3_f097_cond := VAR_uint7_0_0_bit_math_h_l14_c10_592f_return_output;
     VAR_layer1_node0_MUX_bit_math_h_l728_c3_2ff0_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node10_MUX_bit_math_h_l838_c3_cc59_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node11_MUX_bit_math_h_l849_c3_6ba8_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node12_MUX_bit_math_h_l860_c3_e057_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node13_MUX_bit_math_h_l871_c3_aad3_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node14_MUX_bit_math_h_l882_c3_0d3c_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node15_MUX_bit_math_h_l893_c3_6301_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node16_MUX_bit_math_h_l904_c3_60f0_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node17_MUX_bit_math_h_l915_c3_d47f_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node18_MUX_bit_math_h_l926_c3_678f_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node19_MUX_bit_math_h_l937_c3_eb8f_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l739_c3_8d8d_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node20_MUX_bit_math_h_l948_c3_588a_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node21_MUX_bit_math_h_l959_c3_1823_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node22_MUX_bit_math_h_l970_c3_6904_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node23_MUX_bit_math_h_l981_c3_f890_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node24_MUX_bit_math_h_l992_c3_4e65_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node25_MUX_bit_math_h_l1003_c3_f943_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node26_MUX_bit_math_h_l1014_c3_aa20_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node28_MUX_bit_math_h_l1036_c3_85a0_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node29_MUX_bit_math_h_l1047_c3_953f_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l750_c3_7ed6_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node31_MUX_bit_math_h_l1069_c3_82fc_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l761_c3_68af_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node4_MUX_bit_math_h_l772_c3_e8c5_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node5_MUX_bit_math_h_l783_c3_7ab9_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node6_MUX_bit_math_h_l794_c3_1dbe_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node7_MUX_bit_math_h_l805_c3_6dfe_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node8_MUX_bit_math_h_l816_c3_5d19_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer1_node9_MUX_bit_math_h_l827_c3_fe3d_cond := VAR_uint7_1_1_bit_math_h_l724_c10_7c0a_return_output;
     VAR_layer2_node0_MUX_bit_math_h_l1086_c3_4e60_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_12df_return_output;
     VAR_layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_12df_return_output;
     VAR_layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_12df_return_output;
     VAR_layer2_node12_MUX_bit_math_h_l1218_c3_0726_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_12df_return_output;
     VAR_layer2_node13_MUX_bit_math_h_l1229_c3_754d_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_12df_return_output;
     VAR_layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_12df_return_output;
     VAR_layer2_node15_MUX_bit_math_h_l1251_c3_57b2_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_12df_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l1097_c3_12bb_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_12df_return_output;
     VAR_layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_12df_return_output;
     VAR_layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_12df_return_output;
     VAR_layer2_node4_MUX_bit_math_h_l1130_c3_3de0_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_12df_return_output;
     VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_12df_return_output;
     VAR_layer2_node6_MUX_bit_math_h_l1152_c3_3828_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_12df_return_output;
     VAR_layer2_node7_MUX_bit_math_h_l1163_c3_f226_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_12df_return_output;
     VAR_layer2_node8_MUX_bit_math_h_l1174_c3_49b7_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_12df_return_output;
     VAR_layer2_node9_MUX_bit_math_h_l1185_c3_934f_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_12df_return_output;
     VAR_layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_4cf0_return_output;
     VAR_layer3_node1_MUX_bit_math_h_l1279_c3_73ae_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_4cf0_return_output;
     VAR_layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_4cf0_return_output;
     VAR_layer3_node3_MUX_bit_math_h_l1301_c3_827d_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_4cf0_return_output;
     VAR_layer3_node4_MUX_bit_math_h_l1312_c3_ca04_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_4cf0_return_output;
     VAR_layer3_node5_MUX_bit_math_h_l1323_c3_56dd_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_4cf0_return_output;
     VAR_layer3_node6_MUX_bit_math_h_l1334_c3_07bd_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_4cf0_return_output;
     VAR_layer3_node7_MUX_bit_math_h_l1345_c3_5a50_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_4cf0_return_output;
     VAR_layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_cond := VAR_uint7_4_4_bit_math_h_l1358_c10_0af5_return_output;
     VAR_layer4_node1_MUX_bit_math_h_l1373_c3_402b_cond := VAR_uint7_4_4_bit_math_h_l1358_c10_0af5_return_output;
     VAR_layer4_node2_MUX_bit_math_h_l1384_c3_5f80_cond := VAR_uint7_4_4_bit_math_h_l1358_c10_0af5_return_output;
     VAR_layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_cond := VAR_uint7_4_4_bit_math_h_l1358_c10_0af5_return_output;
     VAR_layer5_node0_MUX_bit_math_h_l1412_c3_19e3_cond := VAR_uint7_5_5_bit_math_h_l1408_c10_41c5_return_output;
     VAR_layer5_node1_MUX_bit_math_h_l1423_c3_11f1_cond := VAR_uint7_5_5_bit_math_h_l1408_c10_41c5_return_output;
     VAR_layer6_node0_MUX_bit_math_h_l1440_c3_f906_cond := VAR_uint7_6_6_bit_math_h_l1436_c10_c6df_return_output;
     -- layer0_node14_MUX[bit_math_h_l172_c3_ad25] LATENCY=0
     -- Inputs
     layer0_node14_MUX_bit_math_h_l172_c3_ad25_cond <= VAR_layer0_node14_MUX_bit_math_h_l172_c3_ad25_cond;
     layer0_node14_MUX_bit_math_h_l172_c3_ad25_iftrue <= VAR_layer0_node14_MUX_bit_math_h_l172_c3_ad25_iftrue;
     layer0_node14_MUX_bit_math_h_l172_c3_ad25_iffalse <= VAR_layer0_node14_MUX_bit_math_h_l172_c3_ad25_iffalse;
     -- Outputs
     VAR_layer0_node14_MUX_bit_math_h_l172_c3_ad25_return_output := layer0_node14_MUX_bit_math_h_l172_c3_ad25_return_output;

     -- layer0_node26_MUX[bit_math_h_l304_c3_7f9b] LATENCY=0
     -- Inputs
     layer0_node26_MUX_bit_math_h_l304_c3_7f9b_cond <= VAR_layer0_node26_MUX_bit_math_h_l304_c3_7f9b_cond;
     layer0_node26_MUX_bit_math_h_l304_c3_7f9b_iftrue <= VAR_layer0_node26_MUX_bit_math_h_l304_c3_7f9b_iftrue;
     layer0_node26_MUX_bit_math_h_l304_c3_7f9b_iffalse <= VAR_layer0_node26_MUX_bit_math_h_l304_c3_7f9b_iffalse;
     -- Outputs
     VAR_layer0_node26_MUX_bit_math_h_l304_c3_7f9b_return_output := layer0_node26_MUX_bit_math_h_l304_c3_7f9b_return_output;

     -- layer0_node23_MUX[bit_math_h_l271_c3_86c3] LATENCY=0
     -- Inputs
     layer0_node23_MUX_bit_math_h_l271_c3_86c3_cond <= VAR_layer0_node23_MUX_bit_math_h_l271_c3_86c3_cond;
     layer0_node23_MUX_bit_math_h_l271_c3_86c3_iftrue <= VAR_layer0_node23_MUX_bit_math_h_l271_c3_86c3_iftrue;
     layer0_node23_MUX_bit_math_h_l271_c3_86c3_iffalse <= VAR_layer0_node23_MUX_bit_math_h_l271_c3_86c3_iffalse;
     -- Outputs
     VAR_layer0_node23_MUX_bit_math_h_l271_c3_86c3_return_output := layer0_node23_MUX_bit_math_h_l271_c3_86c3_return_output;

     -- layer0_node42_MUX[bit_math_h_l480_c3_c677] LATENCY=0
     -- Inputs
     layer0_node42_MUX_bit_math_h_l480_c3_c677_cond <= VAR_layer0_node42_MUX_bit_math_h_l480_c3_c677_cond;
     layer0_node42_MUX_bit_math_h_l480_c3_c677_iftrue <= VAR_layer0_node42_MUX_bit_math_h_l480_c3_c677_iftrue;
     layer0_node42_MUX_bit_math_h_l480_c3_c677_iffalse <= VAR_layer0_node42_MUX_bit_math_h_l480_c3_c677_iffalse;
     -- Outputs
     VAR_layer0_node42_MUX_bit_math_h_l480_c3_c677_return_output := layer0_node42_MUX_bit_math_h_l480_c3_c677_return_output;

     -- layer0_node57_MUX[bit_math_h_l645_c3_cec5] LATENCY=0
     -- Inputs
     layer0_node57_MUX_bit_math_h_l645_c3_cec5_cond <= VAR_layer0_node57_MUX_bit_math_h_l645_c3_cec5_cond;
     layer0_node57_MUX_bit_math_h_l645_c3_cec5_iftrue <= VAR_layer0_node57_MUX_bit_math_h_l645_c3_cec5_iftrue;
     layer0_node57_MUX_bit_math_h_l645_c3_cec5_iffalse <= VAR_layer0_node57_MUX_bit_math_h_l645_c3_cec5_iffalse;
     -- Outputs
     VAR_layer0_node57_MUX_bit_math_h_l645_c3_cec5_return_output := layer0_node57_MUX_bit_math_h_l645_c3_cec5_return_output;

     -- layer0_node11_MUX[bit_math_h_l139_c3_3ab9] LATENCY=0
     -- Inputs
     layer0_node11_MUX_bit_math_h_l139_c3_3ab9_cond <= VAR_layer0_node11_MUX_bit_math_h_l139_c3_3ab9_cond;
     layer0_node11_MUX_bit_math_h_l139_c3_3ab9_iftrue <= VAR_layer0_node11_MUX_bit_math_h_l139_c3_3ab9_iftrue;
     layer0_node11_MUX_bit_math_h_l139_c3_3ab9_iffalse <= VAR_layer0_node11_MUX_bit_math_h_l139_c3_3ab9_iffalse;
     -- Outputs
     VAR_layer0_node11_MUX_bit_math_h_l139_c3_3ab9_return_output := layer0_node11_MUX_bit_math_h_l139_c3_3ab9_return_output;

     -- layer0_node16_MUX[bit_math_h_l194_c3_5393] LATENCY=0
     -- Inputs
     layer0_node16_MUX_bit_math_h_l194_c3_5393_cond <= VAR_layer0_node16_MUX_bit_math_h_l194_c3_5393_cond;
     layer0_node16_MUX_bit_math_h_l194_c3_5393_iftrue <= VAR_layer0_node16_MUX_bit_math_h_l194_c3_5393_iftrue;
     layer0_node16_MUX_bit_math_h_l194_c3_5393_iffalse <= VAR_layer0_node16_MUX_bit_math_h_l194_c3_5393_iffalse;
     -- Outputs
     VAR_layer0_node16_MUX_bit_math_h_l194_c3_5393_return_output := layer0_node16_MUX_bit_math_h_l194_c3_5393_return_output;

     -- layer0_node5_MUX[bit_math_h_l73_c3_282b] LATENCY=0
     -- Inputs
     layer0_node5_MUX_bit_math_h_l73_c3_282b_cond <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_282b_cond;
     layer0_node5_MUX_bit_math_h_l73_c3_282b_iftrue <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_282b_iftrue;
     layer0_node5_MUX_bit_math_h_l73_c3_282b_iffalse <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_282b_iffalse;
     -- Outputs
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_282b_return_output := layer0_node5_MUX_bit_math_h_l73_c3_282b_return_output;

     -- layer0_node0_MUX[bit_math_h_l18_c3_5c06] LATENCY=0
     -- Inputs
     layer0_node0_MUX_bit_math_h_l18_c3_5c06_cond <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_5c06_cond;
     layer0_node0_MUX_bit_math_h_l18_c3_5c06_iftrue <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_5c06_iftrue;
     layer0_node0_MUX_bit_math_h_l18_c3_5c06_iffalse <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_5c06_iffalse;
     -- Outputs
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_5c06_return_output := layer0_node0_MUX_bit_math_h_l18_c3_5c06_return_output;

     -- layer0_node36_MUX[bit_math_h_l414_c3_cd2c] LATENCY=0
     -- Inputs
     layer0_node36_MUX_bit_math_h_l414_c3_cd2c_cond <= VAR_layer0_node36_MUX_bit_math_h_l414_c3_cd2c_cond;
     layer0_node36_MUX_bit_math_h_l414_c3_cd2c_iftrue <= VAR_layer0_node36_MUX_bit_math_h_l414_c3_cd2c_iftrue;
     layer0_node36_MUX_bit_math_h_l414_c3_cd2c_iffalse <= VAR_layer0_node36_MUX_bit_math_h_l414_c3_cd2c_iffalse;
     -- Outputs
     VAR_layer0_node36_MUX_bit_math_h_l414_c3_cd2c_return_output := layer0_node36_MUX_bit_math_h_l414_c3_cd2c_return_output;

     -- layer0_node7_MUX[bit_math_h_l95_c3_567b] LATENCY=0
     -- Inputs
     layer0_node7_MUX_bit_math_h_l95_c3_567b_cond <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_567b_cond;
     layer0_node7_MUX_bit_math_h_l95_c3_567b_iftrue <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_567b_iftrue;
     layer0_node7_MUX_bit_math_h_l95_c3_567b_iffalse <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_567b_iffalse;
     -- Outputs
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_567b_return_output := layer0_node7_MUX_bit_math_h_l95_c3_567b_return_output;

     -- layer0_node59_MUX[bit_math_h_l667_c3_672d] LATENCY=0
     -- Inputs
     layer0_node59_MUX_bit_math_h_l667_c3_672d_cond <= VAR_layer0_node59_MUX_bit_math_h_l667_c3_672d_cond;
     layer0_node59_MUX_bit_math_h_l667_c3_672d_iftrue <= VAR_layer0_node59_MUX_bit_math_h_l667_c3_672d_iftrue;
     layer0_node59_MUX_bit_math_h_l667_c3_672d_iffalse <= VAR_layer0_node59_MUX_bit_math_h_l667_c3_672d_iffalse;
     -- Outputs
     VAR_layer0_node59_MUX_bit_math_h_l667_c3_672d_return_output := layer0_node59_MUX_bit_math_h_l667_c3_672d_return_output;

     -- layer0_node6_MUX[bit_math_h_l84_c3_62f1] LATENCY=0
     -- Inputs
     layer0_node6_MUX_bit_math_h_l84_c3_62f1_cond <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_62f1_cond;
     layer0_node6_MUX_bit_math_h_l84_c3_62f1_iftrue <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_62f1_iftrue;
     layer0_node6_MUX_bit_math_h_l84_c3_62f1_iffalse <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_62f1_iffalse;
     -- Outputs
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_62f1_return_output := layer0_node6_MUX_bit_math_h_l84_c3_62f1_return_output;

     -- layer0_node28_MUX[bit_math_h_l326_c3_12a3] LATENCY=0
     -- Inputs
     layer0_node28_MUX_bit_math_h_l326_c3_12a3_cond <= VAR_layer0_node28_MUX_bit_math_h_l326_c3_12a3_cond;
     layer0_node28_MUX_bit_math_h_l326_c3_12a3_iftrue <= VAR_layer0_node28_MUX_bit_math_h_l326_c3_12a3_iftrue;
     layer0_node28_MUX_bit_math_h_l326_c3_12a3_iffalse <= VAR_layer0_node28_MUX_bit_math_h_l326_c3_12a3_iffalse;
     -- Outputs
     VAR_layer0_node28_MUX_bit_math_h_l326_c3_12a3_return_output := layer0_node28_MUX_bit_math_h_l326_c3_12a3_return_output;

     -- layer0_node45_MUX[bit_math_h_l513_c3_b86e] LATENCY=0
     -- Inputs
     layer0_node45_MUX_bit_math_h_l513_c3_b86e_cond <= VAR_layer0_node45_MUX_bit_math_h_l513_c3_b86e_cond;
     layer0_node45_MUX_bit_math_h_l513_c3_b86e_iftrue <= VAR_layer0_node45_MUX_bit_math_h_l513_c3_b86e_iftrue;
     layer0_node45_MUX_bit_math_h_l513_c3_b86e_iffalse <= VAR_layer0_node45_MUX_bit_math_h_l513_c3_b86e_iffalse;
     -- Outputs
     VAR_layer0_node45_MUX_bit_math_h_l513_c3_b86e_return_output := layer0_node45_MUX_bit_math_h_l513_c3_b86e_return_output;

     -- layer0_node22_MUX[bit_math_h_l260_c3_321e] LATENCY=0
     -- Inputs
     layer0_node22_MUX_bit_math_h_l260_c3_321e_cond <= VAR_layer0_node22_MUX_bit_math_h_l260_c3_321e_cond;
     layer0_node22_MUX_bit_math_h_l260_c3_321e_iftrue <= VAR_layer0_node22_MUX_bit_math_h_l260_c3_321e_iftrue;
     layer0_node22_MUX_bit_math_h_l260_c3_321e_iffalse <= VAR_layer0_node22_MUX_bit_math_h_l260_c3_321e_iffalse;
     -- Outputs
     VAR_layer0_node22_MUX_bit_math_h_l260_c3_321e_return_output := layer0_node22_MUX_bit_math_h_l260_c3_321e_return_output;

     -- layer0_node61_MUX[bit_math_h_l689_c3_be95] LATENCY=0
     -- Inputs
     layer0_node61_MUX_bit_math_h_l689_c3_be95_cond <= VAR_layer0_node61_MUX_bit_math_h_l689_c3_be95_cond;
     layer0_node61_MUX_bit_math_h_l689_c3_be95_iftrue <= VAR_layer0_node61_MUX_bit_math_h_l689_c3_be95_iftrue;
     layer0_node61_MUX_bit_math_h_l689_c3_be95_iffalse <= VAR_layer0_node61_MUX_bit_math_h_l689_c3_be95_iffalse;
     -- Outputs
     VAR_layer0_node61_MUX_bit_math_h_l689_c3_be95_return_output := layer0_node61_MUX_bit_math_h_l689_c3_be95_return_output;

     -- layer0_node30_MUX[bit_math_h_l348_c3_8c5c] LATENCY=0
     -- Inputs
     layer0_node30_MUX_bit_math_h_l348_c3_8c5c_cond <= VAR_layer0_node30_MUX_bit_math_h_l348_c3_8c5c_cond;
     layer0_node30_MUX_bit_math_h_l348_c3_8c5c_iftrue <= VAR_layer0_node30_MUX_bit_math_h_l348_c3_8c5c_iftrue;
     layer0_node30_MUX_bit_math_h_l348_c3_8c5c_iffalse <= VAR_layer0_node30_MUX_bit_math_h_l348_c3_8c5c_iffalse;
     -- Outputs
     VAR_layer0_node30_MUX_bit_math_h_l348_c3_8c5c_return_output := layer0_node30_MUX_bit_math_h_l348_c3_8c5c_return_output;

     -- layer0_node31_MUX[bit_math_h_l359_c3_d6b9] LATENCY=0
     -- Inputs
     layer0_node31_MUX_bit_math_h_l359_c3_d6b9_cond <= VAR_layer0_node31_MUX_bit_math_h_l359_c3_d6b9_cond;
     layer0_node31_MUX_bit_math_h_l359_c3_d6b9_iftrue <= VAR_layer0_node31_MUX_bit_math_h_l359_c3_d6b9_iftrue;
     layer0_node31_MUX_bit_math_h_l359_c3_d6b9_iffalse <= VAR_layer0_node31_MUX_bit_math_h_l359_c3_d6b9_iffalse;
     -- Outputs
     VAR_layer0_node31_MUX_bit_math_h_l359_c3_d6b9_return_output := layer0_node31_MUX_bit_math_h_l359_c3_d6b9_return_output;

     -- layer0_node35_MUX[bit_math_h_l403_c3_683e] LATENCY=0
     -- Inputs
     layer0_node35_MUX_bit_math_h_l403_c3_683e_cond <= VAR_layer0_node35_MUX_bit_math_h_l403_c3_683e_cond;
     layer0_node35_MUX_bit_math_h_l403_c3_683e_iftrue <= VAR_layer0_node35_MUX_bit_math_h_l403_c3_683e_iftrue;
     layer0_node35_MUX_bit_math_h_l403_c3_683e_iffalse <= VAR_layer0_node35_MUX_bit_math_h_l403_c3_683e_iffalse;
     -- Outputs
     VAR_layer0_node35_MUX_bit_math_h_l403_c3_683e_return_output := layer0_node35_MUX_bit_math_h_l403_c3_683e_return_output;

     -- layer0_node21_MUX[bit_math_h_l249_c3_8f8c] LATENCY=0
     -- Inputs
     layer0_node21_MUX_bit_math_h_l249_c3_8f8c_cond <= VAR_layer0_node21_MUX_bit_math_h_l249_c3_8f8c_cond;
     layer0_node21_MUX_bit_math_h_l249_c3_8f8c_iftrue <= VAR_layer0_node21_MUX_bit_math_h_l249_c3_8f8c_iftrue;
     layer0_node21_MUX_bit_math_h_l249_c3_8f8c_iffalse <= VAR_layer0_node21_MUX_bit_math_h_l249_c3_8f8c_iffalse;
     -- Outputs
     VAR_layer0_node21_MUX_bit_math_h_l249_c3_8f8c_return_output := layer0_node21_MUX_bit_math_h_l249_c3_8f8c_return_output;

     -- layer0_node58_MUX[bit_math_h_l656_c3_312b] LATENCY=0
     -- Inputs
     layer0_node58_MUX_bit_math_h_l656_c3_312b_cond <= VAR_layer0_node58_MUX_bit_math_h_l656_c3_312b_cond;
     layer0_node58_MUX_bit_math_h_l656_c3_312b_iftrue <= VAR_layer0_node58_MUX_bit_math_h_l656_c3_312b_iftrue;
     layer0_node58_MUX_bit_math_h_l656_c3_312b_iffalse <= VAR_layer0_node58_MUX_bit_math_h_l656_c3_312b_iffalse;
     -- Outputs
     VAR_layer0_node58_MUX_bit_math_h_l656_c3_312b_return_output := layer0_node58_MUX_bit_math_h_l656_c3_312b_return_output;

     -- layer0_node63_MUX[bit_math_h_l711_c3_45fc] LATENCY=0
     -- Inputs
     layer0_node63_MUX_bit_math_h_l711_c3_45fc_cond <= VAR_layer0_node63_MUX_bit_math_h_l711_c3_45fc_cond;
     layer0_node63_MUX_bit_math_h_l711_c3_45fc_iftrue <= VAR_layer0_node63_MUX_bit_math_h_l711_c3_45fc_iftrue;
     layer0_node63_MUX_bit_math_h_l711_c3_45fc_iffalse <= VAR_layer0_node63_MUX_bit_math_h_l711_c3_45fc_iffalse;
     -- Outputs
     VAR_layer0_node63_MUX_bit_math_h_l711_c3_45fc_return_output := layer0_node63_MUX_bit_math_h_l711_c3_45fc_return_output;

     -- layer0_node54_MUX[bit_math_h_l612_c3_cab9] LATENCY=0
     -- Inputs
     layer0_node54_MUX_bit_math_h_l612_c3_cab9_cond <= VAR_layer0_node54_MUX_bit_math_h_l612_c3_cab9_cond;
     layer0_node54_MUX_bit_math_h_l612_c3_cab9_iftrue <= VAR_layer0_node54_MUX_bit_math_h_l612_c3_cab9_iftrue;
     layer0_node54_MUX_bit_math_h_l612_c3_cab9_iffalse <= VAR_layer0_node54_MUX_bit_math_h_l612_c3_cab9_iffalse;
     -- Outputs
     VAR_layer0_node54_MUX_bit_math_h_l612_c3_cab9_return_output := layer0_node54_MUX_bit_math_h_l612_c3_cab9_return_output;

     -- layer0_node15_MUX[bit_math_h_l183_c3_dacd] LATENCY=0
     -- Inputs
     layer0_node15_MUX_bit_math_h_l183_c3_dacd_cond <= VAR_layer0_node15_MUX_bit_math_h_l183_c3_dacd_cond;
     layer0_node15_MUX_bit_math_h_l183_c3_dacd_iftrue <= VAR_layer0_node15_MUX_bit_math_h_l183_c3_dacd_iftrue;
     layer0_node15_MUX_bit_math_h_l183_c3_dacd_iffalse <= VAR_layer0_node15_MUX_bit_math_h_l183_c3_dacd_iffalse;
     -- Outputs
     VAR_layer0_node15_MUX_bit_math_h_l183_c3_dacd_return_output := layer0_node15_MUX_bit_math_h_l183_c3_dacd_return_output;

     -- layer0_node10_MUX[bit_math_h_l128_c3_0e6c] LATENCY=0
     -- Inputs
     layer0_node10_MUX_bit_math_h_l128_c3_0e6c_cond <= VAR_layer0_node10_MUX_bit_math_h_l128_c3_0e6c_cond;
     layer0_node10_MUX_bit_math_h_l128_c3_0e6c_iftrue <= VAR_layer0_node10_MUX_bit_math_h_l128_c3_0e6c_iftrue;
     layer0_node10_MUX_bit_math_h_l128_c3_0e6c_iffalse <= VAR_layer0_node10_MUX_bit_math_h_l128_c3_0e6c_iffalse;
     -- Outputs
     VAR_layer0_node10_MUX_bit_math_h_l128_c3_0e6c_return_output := layer0_node10_MUX_bit_math_h_l128_c3_0e6c_return_output;

     -- layer0_node1_MUX[bit_math_h_l29_c3_fa46] LATENCY=0
     -- Inputs
     layer0_node1_MUX_bit_math_h_l29_c3_fa46_cond <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_fa46_cond;
     layer0_node1_MUX_bit_math_h_l29_c3_fa46_iftrue <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_fa46_iftrue;
     layer0_node1_MUX_bit_math_h_l29_c3_fa46_iffalse <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_fa46_iffalse;
     -- Outputs
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_fa46_return_output := layer0_node1_MUX_bit_math_h_l29_c3_fa46_return_output;

     -- layer0_node44_MUX[bit_math_h_l502_c3_6b96] LATENCY=0
     -- Inputs
     layer0_node44_MUX_bit_math_h_l502_c3_6b96_cond <= VAR_layer0_node44_MUX_bit_math_h_l502_c3_6b96_cond;
     layer0_node44_MUX_bit_math_h_l502_c3_6b96_iftrue <= VAR_layer0_node44_MUX_bit_math_h_l502_c3_6b96_iftrue;
     layer0_node44_MUX_bit_math_h_l502_c3_6b96_iffalse <= VAR_layer0_node44_MUX_bit_math_h_l502_c3_6b96_iffalse;
     -- Outputs
     VAR_layer0_node44_MUX_bit_math_h_l502_c3_6b96_return_output := layer0_node44_MUX_bit_math_h_l502_c3_6b96_return_output;

     -- layer0_node8_MUX[bit_math_h_l106_c3_47e5] LATENCY=0
     -- Inputs
     layer0_node8_MUX_bit_math_h_l106_c3_47e5_cond <= VAR_layer0_node8_MUX_bit_math_h_l106_c3_47e5_cond;
     layer0_node8_MUX_bit_math_h_l106_c3_47e5_iftrue <= VAR_layer0_node8_MUX_bit_math_h_l106_c3_47e5_iftrue;
     layer0_node8_MUX_bit_math_h_l106_c3_47e5_iffalse <= VAR_layer0_node8_MUX_bit_math_h_l106_c3_47e5_iffalse;
     -- Outputs
     VAR_layer0_node8_MUX_bit_math_h_l106_c3_47e5_return_output := layer0_node8_MUX_bit_math_h_l106_c3_47e5_return_output;

     -- layer0_node34_MUX[bit_math_h_l392_c3_f617] LATENCY=0
     -- Inputs
     layer0_node34_MUX_bit_math_h_l392_c3_f617_cond <= VAR_layer0_node34_MUX_bit_math_h_l392_c3_f617_cond;
     layer0_node34_MUX_bit_math_h_l392_c3_f617_iftrue <= VAR_layer0_node34_MUX_bit_math_h_l392_c3_f617_iftrue;
     layer0_node34_MUX_bit_math_h_l392_c3_f617_iffalse <= VAR_layer0_node34_MUX_bit_math_h_l392_c3_f617_iffalse;
     -- Outputs
     VAR_layer0_node34_MUX_bit_math_h_l392_c3_f617_return_output := layer0_node34_MUX_bit_math_h_l392_c3_f617_return_output;

     -- layer0_node49_MUX[bit_math_h_l557_c3_3410] LATENCY=0
     -- Inputs
     layer0_node49_MUX_bit_math_h_l557_c3_3410_cond <= VAR_layer0_node49_MUX_bit_math_h_l557_c3_3410_cond;
     layer0_node49_MUX_bit_math_h_l557_c3_3410_iftrue <= VAR_layer0_node49_MUX_bit_math_h_l557_c3_3410_iftrue;
     layer0_node49_MUX_bit_math_h_l557_c3_3410_iffalse <= VAR_layer0_node49_MUX_bit_math_h_l557_c3_3410_iffalse;
     -- Outputs
     VAR_layer0_node49_MUX_bit_math_h_l557_c3_3410_return_output := layer0_node49_MUX_bit_math_h_l557_c3_3410_return_output;

     -- layer0_node43_MUX[bit_math_h_l491_c3_2838] LATENCY=0
     -- Inputs
     layer0_node43_MUX_bit_math_h_l491_c3_2838_cond <= VAR_layer0_node43_MUX_bit_math_h_l491_c3_2838_cond;
     layer0_node43_MUX_bit_math_h_l491_c3_2838_iftrue <= VAR_layer0_node43_MUX_bit_math_h_l491_c3_2838_iftrue;
     layer0_node43_MUX_bit_math_h_l491_c3_2838_iffalse <= VAR_layer0_node43_MUX_bit_math_h_l491_c3_2838_iffalse;
     -- Outputs
     VAR_layer0_node43_MUX_bit_math_h_l491_c3_2838_return_output := layer0_node43_MUX_bit_math_h_l491_c3_2838_return_output;

     -- layer0_node55_MUX[bit_math_h_l623_c3_2e5e] LATENCY=0
     -- Inputs
     layer0_node55_MUX_bit_math_h_l623_c3_2e5e_cond <= VAR_layer0_node55_MUX_bit_math_h_l623_c3_2e5e_cond;
     layer0_node55_MUX_bit_math_h_l623_c3_2e5e_iftrue <= VAR_layer0_node55_MUX_bit_math_h_l623_c3_2e5e_iftrue;
     layer0_node55_MUX_bit_math_h_l623_c3_2e5e_iffalse <= VAR_layer0_node55_MUX_bit_math_h_l623_c3_2e5e_iffalse;
     -- Outputs
     VAR_layer0_node55_MUX_bit_math_h_l623_c3_2e5e_return_output := layer0_node55_MUX_bit_math_h_l623_c3_2e5e_return_output;

     -- layer0_node51_MUX[bit_math_h_l579_c3_8398] LATENCY=0
     -- Inputs
     layer0_node51_MUX_bit_math_h_l579_c3_8398_cond <= VAR_layer0_node51_MUX_bit_math_h_l579_c3_8398_cond;
     layer0_node51_MUX_bit_math_h_l579_c3_8398_iftrue <= VAR_layer0_node51_MUX_bit_math_h_l579_c3_8398_iftrue;
     layer0_node51_MUX_bit_math_h_l579_c3_8398_iffalse <= VAR_layer0_node51_MUX_bit_math_h_l579_c3_8398_iffalse;
     -- Outputs
     VAR_layer0_node51_MUX_bit_math_h_l579_c3_8398_return_output := layer0_node51_MUX_bit_math_h_l579_c3_8398_return_output;

     -- layer0_node52_MUX[bit_math_h_l590_c3_6d3d] LATENCY=0
     -- Inputs
     layer0_node52_MUX_bit_math_h_l590_c3_6d3d_cond <= VAR_layer0_node52_MUX_bit_math_h_l590_c3_6d3d_cond;
     layer0_node52_MUX_bit_math_h_l590_c3_6d3d_iftrue <= VAR_layer0_node52_MUX_bit_math_h_l590_c3_6d3d_iftrue;
     layer0_node52_MUX_bit_math_h_l590_c3_6d3d_iffalse <= VAR_layer0_node52_MUX_bit_math_h_l590_c3_6d3d_iffalse;
     -- Outputs
     VAR_layer0_node52_MUX_bit_math_h_l590_c3_6d3d_return_output := layer0_node52_MUX_bit_math_h_l590_c3_6d3d_return_output;

     -- layer0_node19_MUX[bit_math_h_l227_c3_1dae] LATENCY=0
     -- Inputs
     layer0_node19_MUX_bit_math_h_l227_c3_1dae_cond <= VAR_layer0_node19_MUX_bit_math_h_l227_c3_1dae_cond;
     layer0_node19_MUX_bit_math_h_l227_c3_1dae_iftrue <= VAR_layer0_node19_MUX_bit_math_h_l227_c3_1dae_iftrue;
     layer0_node19_MUX_bit_math_h_l227_c3_1dae_iffalse <= VAR_layer0_node19_MUX_bit_math_h_l227_c3_1dae_iffalse;
     -- Outputs
     VAR_layer0_node19_MUX_bit_math_h_l227_c3_1dae_return_output := layer0_node19_MUX_bit_math_h_l227_c3_1dae_return_output;

     -- layer0_node9_MUX[bit_math_h_l117_c3_f097] LATENCY=0
     -- Inputs
     layer0_node9_MUX_bit_math_h_l117_c3_f097_cond <= VAR_layer0_node9_MUX_bit_math_h_l117_c3_f097_cond;
     layer0_node9_MUX_bit_math_h_l117_c3_f097_iftrue <= VAR_layer0_node9_MUX_bit_math_h_l117_c3_f097_iftrue;
     layer0_node9_MUX_bit_math_h_l117_c3_f097_iffalse <= VAR_layer0_node9_MUX_bit_math_h_l117_c3_f097_iffalse;
     -- Outputs
     VAR_layer0_node9_MUX_bit_math_h_l117_c3_f097_return_output := layer0_node9_MUX_bit_math_h_l117_c3_f097_return_output;

     -- layer0_node2_MUX[bit_math_h_l40_c3_f68a] LATENCY=0
     -- Inputs
     layer0_node2_MUX_bit_math_h_l40_c3_f68a_cond <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_f68a_cond;
     layer0_node2_MUX_bit_math_h_l40_c3_f68a_iftrue <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_f68a_iftrue;
     layer0_node2_MUX_bit_math_h_l40_c3_f68a_iffalse <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_f68a_iffalse;
     -- Outputs
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_f68a_return_output := layer0_node2_MUX_bit_math_h_l40_c3_f68a_return_output;

     -- layer0_node12_MUX[bit_math_h_l150_c3_e611] LATENCY=0
     -- Inputs
     layer0_node12_MUX_bit_math_h_l150_c3_e611_cond <= VAR_layer0_node12_MUX_bit_math_h_l150_c3_e611_cond;
     layer0_node12_MUX_bit_math_h_l150_c3_e611_iftrue <= VAR_layer0_node12_MUX_bit_math_h_l150_c3_e611_iftrue;
     layer0_node12_MUX_bit_math_h_l150_c3_e611_iffalse <= VAR_layer0_node12_MUX_bit_math_h_l150_c3_e611_iffalse;
     -- Outputs
     VAR_layer0_node12_MUX_bit_math_h_l150_c3_e611_return_output := layer0_node12_MUX_bit_math_h_l150_c3_e611_return_output;

     -- layer0_node41_MUX[bit_math_h_l469_c3_b3bf] LATENCY=0
     -- Inputs
     layer0_node41_MUX_bit_math_h_l469_c3_b3bf_cond <= VAR_layer0_node41_MUX_bit_math_h_l469_c3_b3bf_cond;
     layer0_node41_MUX_bit_math_h_l469_c3_b3bf_iftrue <= VAR_layer0_node41_MUX_bit_math_h_l469_c3_b3bf_iftrue;
     layer0_node41_MUX_bit_math_h_l469_c3_b3bf_iffalse <= VAR_layer0_node41_MUX_bit_math_h_l469_c3_b3bf_iffalse;
     -- Outputs
     VAR_layer0_node41_MUX_bit_math_h_l469_c3_b3bf_return_output := layer0_node41_MUX_bit_math_h_l469_c3_b3bf_return_output;

     -- layer0_node17_MUX[bit_math_h_l205_c3_4246] LATENCY=0
     -- Inputs
     layer0_node17_MUX_bit_math_h_l205_c3_4246_cond <= VAR_layer0_node17_MUX_bit_math_h_l205_c3_4246_cond;
     layer0_node17_MUX_bit_math_h_l205_c3_4246_iftrue <= VAR_layer0_node17_MUX_bit_math_h_l205_c3_4246_iftrue;
     layer0_node17_MUX_bit_math_h_l205_c3_4246_iffalse <= VAR_layer0_node17_MUX_bit_math_h_l205_c3_4246_iffalse;
     -- Outputs
     VAR_layer0_node17_MUX_bit_math_h_l205_c3_4246_return_output := layer0_node17_MUX_bit_math_h_l205_c3_4246_return_output;

     -- layer0_node48_MUX[bit_math_h_l546_c3_5be4] LATENCY=0
     -- Inputs
     layer0_node48_MUX_bit_math_h_l546_c3_5be4_cond <= VAR_layer0_node48_MUX_bit_math_h_l546_c3_5be4_cond;
     layer0_node48_MUX_bit_math_h_l546_c3_5be4_iftrue <= VAR_layer0_node48_MUX_bit_math_h_l546_c3_5be4_iftrue;
     layer0_node48_MUX_bit_math_h_l546_c3_5be4_iffalse <= VAR_layer0_node48_MUX_bit_math_h_l546_c3_5be4_iffalse;
     -- Outputs
     VAR_layer0_node48_MUX_bit_math_h_l546_c3_5be4_return_output := layer0_node48_MUX_bit_math_h_l546_c3_5be4_return_output;

     -- layer0_node25_MUX[bit_math_h_l293_c3_ece2] LATENCY=0
     -- Inputs
     layer0_node25_MUX_bit_math_h_l293_c3_ece2_cond <= VAR_layer0_node25_MUX_bit_math_h_l293_c3_ece2_cond;
     layer0_node25_MUX_bit_math_h_l293_c3_ece2_iftrue <= VAR_layer0_node25_MUX_bit_math_h_l293_c3_ece2_iftrue;
     layer0_node25_MUX_bit_math_h_l293_c3_ece2_iffalse <= VAR_layer0_node25_MUX_bit_math_h_l293_c3_ece2_iffalse;
     -- Outputs
     VAR_layer0_node25_MUX_bit_math_h_l293_c3_ece2_return_output := layer0_node25_MUX_bit_math_h_l293_c3_ece2_return_output;

     -- layer0_node4_MUX[bit_math_h_l62_c3_07e7] LATENCY=0
     -- Inputs
     layer0_node4_MUX_bit_math_h_l62_c3_07e7_cond <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_07e7_cond;
     layer0_node4_MUX_bit_math_h_l62_c3_07e7_iftrue <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_07e7_iftrue;
     layer0_node4_MUX_bit_math_h_l62_c3_07e7_iffalse <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_07e7_iffalse;
     -- Outputs
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_07e7_return_output := layer0_node4_MUX_bit_math_h_l62_c3_07e7_return_output;

     -- layer0_node20_MUX[bit_math_h_l238_c3_e7c7] LATENCY=0
     -- Inputs
     layer0_node20_MUX_bit_math_h_l238_c3_e7c7_cond <= VAR_layer0_node20_MUX_bit_math_h_l238_c3_e7c7_cond;
     layer0_node20_MUX_bit_math_h_l238_c3_e7c7_iftrue <= VAR_layer0_node20_MUX_bit_math_h_l238_c3_e7c7_iftrue;
     layer0_node20_MUX_bit_math_h_l238_c3_e7c7_iffalse <= VAR_layer0_node20_MUX_bit_math_h_l238_c3_e7c7_iffalse;
     -- Outputs
     VAR_layer0_node20_MUX_bit_math_h_l238_c3_e7c7_return_output := layer0_node20_MUX_bit_math_h_l238_c3_e7c7_return_output;

     -- layer0_node47_MUX[bit_math_h_l535_c3_21f3] LATENCY=0
     -- Inputs
     layer0_node47_MUX_bit_math_h_l535_c3_21f3_cond <= VAR_layer0_node47_MUX_bit_math_h_l535_c3_21f3_cond;
     layer0_node47_MUX_bit_math_h_l535_c3_21f3_iftrue <= VAR_layer0_node47_MUX_bit_math_h_l535_c3_21f3_iftrue;
     layer0_node47_MUX_bit_math_h_l535_c3_21f3_iffalse <= VAR_layer0_node47_MUX_bit_math_h_l535_c3_21f3_iffalse;
     -- Outputs
     VAR_layer0_node47_MUX_bit_math_h_l535_c3_21f3_return_output := layer0_node47_MUX_bit_math_h_l535_c3_21f3_return_output;

     -- layer0_node62_MUX[bit_math_h_l700_c3_8a98] LATENCY=0
     -- Inputs
     layer0_node62_MUX_bit_math_h_l700_c3_8a98_cond <= VAR_layer0_node62_MUX_bit_math_h_l700_c3_8a98_cond;
     layer0_node62_MUX_bit_math_h_l700_c3_8a98_iftrue <= VAR_layer0_node62_MUX_bit_math_h_l700_c3_8a98_iftrue;
     layer0_node62_MUX_bit_math_h_l700_c3_8a98_iffalse <= VAR_layer0_node62_MUX_bit_math_h_l700_c3_8a98_iffalse;
     -- Outputs
     VAR_layer0_node62_MUX_bit_math_h_l700_c3_8a98_return_output := layer0_node62_MUX_bit_math_h_l700_c3_8a98_return_output;

     -- layer0_node33_MUX[bit_math_h_l381_c3_bdd0] LATENCY=0
     -- Inputs
     layer0_node33_MUX_bit_math_h_l381_c3_bdd0_cond <= VAR_layer0_node33_MUX_bit_math_h_l381_c3_bdd0_cond;
     layer0_node33_MUX_bit_math_h_l381_c3_bdd0_iftrue <= VAR_layer0_node33_MUX_bit_math_h_l381_c3_bdd0_iftrue;
     layer0_node33_MUX_bit_math_h_l381_c3_bdd0_iffalse <= VAR_layer0_node33_MUX_bit_math_h_l381_c3_bdd0_iffalse;
     -- Outputs
     VAR_layer0_node33_MUX_bit_math_h_l381_c3_bdd0_return_output := layer0_node33_MUX_bit_math_h_l381_c3_bdd0_return_output;

     -- layer0_node39_MUX[bit_math_h_l447_c3_b150] LATENCY=0
     -- Inputs
     layer0_node39_MUX_bit_math_h_l447_c3_b150_cond <= VAR_layer0_node39_MUX_bit_math_h_l447_c3_b150_cond;
     layer0_node39_MUX_bit_math_h_l447_c3_b150_iftrue <= VAR_layer0_node39_MUX_bit_math_h_l447_c3_b150_iftrue;
     layer0_node39_MUX_bit_math_h_l447_c3_b150_iffalse <= VAR_layer0_node39_MUX_bit_math_h_l447_c3_b150_iffalse;
     -- Outputs
     VAR_layer0_node39_MUX_bit_math_h_l447_c3_b150_return_output := layer0_node39_MUX_bit_math_h_l447_c3_b150_return_output;

     -- layer0_node13_MUX[bit_math_h_l161_c3_e037] LATENCY=0
     -- Inputs
     layer0_node13_MUX_bit_math_h_l161_c3_e037_cond <= VAR_layer0_node13_MUX_bit_math_h_l161_c3_e037_cond;
     layer0_node13_MUX_bit_math_h_l161_c3_e037_iftrue <= VAR_layer0_node13_MUX_bit_math_h_l161_c3_e037_iftrue;
     layer0_node13_MUX_bit_math_h_l161_c3_e037_iffalse <= VAR_layer0_node13_MUX_bit_math_h_l161_c3_e037_iffalse;
     -- Outputs
     VAR_layer0_node13_MUX_bit_math_h_l161_c3_e037_return_output := layer0_node13_MUX_bit_math_h_l161_c3_e037_return_output;

     -- layer0_node24_MUX[bit_math_h_l282_c3_2992] LATENCY=0
     -- Inputs
     layer0_node24_MUX_bit_math_h_l282_c3_2992_cond <= VAR_layer0_node24_MUX_bit_math_h_l282_c3_2992_cond;
     layer0_node24_MUX_bit_math_h_l282_c3_2992_iftrue <= VAR_layer0_node24_MUX_bit_math_h_l282_c3_2992_iftrue;
     layer0_node24_MUX_bit_math_h_l282_c3_2992_iffalse <= VAR_layer0_node24_MUX_bit_math_h_l282_c3_2992_iffalse;
     -- Outputs
     VAR_layer0_node24_MUX_bit_math_h_l282_c3_2992_return_output := layer0_node24_MUX_bit_math_h_l282_c3_2992_return_output;

     -- layer0_node38_MUX[bit_math_h_l436_c3_c940] LATENCY=0
     -- Inputs
     layer0_node38_MUX_bit_math_h_l436_c3_c940_cond <= VAR_layer0_node38_MUX_bit_math_h_l436_c3_c940_cond;
     layer0_node38_MUX_bit_math_h_l436_c3_c940_iftrue <= VAR_layer0_node38_MUX_bit_math_h_l436_c3_c940_iftrue;
     layer0_node38_MUX_bit_math_h_l436_c3_c940_iffalse <= VAR_layer0_node38_MUX_bit_math_h_l436_c3_c940_iffalse;
     -- Outputs
     VAR_layer0_node38_MUX_bit_math_h_l436_c3_c940_return_output := layer0_node38_MUX_bit_math_h_l436_c3_c940_return_output;

     -- layer0_node60_MUX[bit_math_h_l678_c3_9a42] LATENCY=0
     -- Inputs
     layer0_node60_MUX_bit_math_h_l678_c3_9a42_cond <= VAR_layer0_node60_MUX_bit_math_h_l678_c3_9a42_cond;
     layer0_node60_MUX_bit_math_h_l678_c3_9a42_iftrue <= VAR_layer0_node60_MUX_bit_math_h_l678_c3_9a42_iftrue;
     layer0_node60_MUX_bit_math_h_l678_c3_9a42_iffalse <= VAR_layer0_node60_MUX_bit_math_h_l678_c3_9a42_iffalse;
     -- Outputs
     VAR_layer0_node60_MUX_bit_math_h_l678_c3_9a42_return_output := layer0_node60_MUX_bit_math_h_l678_c3_9a42_return_output;

     -- layer0_node18_MUX[bit_math_h_l216_c3_2748] LATENCY=0
     -- Inputs
     layer0_node18_MUX_bit_math_h_l216_c3_2748_cond <= VAR_layer0_node18_MUX_bit_math_h_l216_c3_2748_cond;
     layer0_node18_MUX_bit_math_h_l216_c3_2748_iftrue <= VAR_layer0_node18_MUX_bit_math_h_l216_c3_2748_iftrue;
     layer0_node18_MUX_bit_math_h_l216_c3_2748_iffalse <= VAR_layer0_node18_MUX_bit_math_h_l216_c3_2748_iffalse;
     -- Outputs
     VAR_layer0_node18_MUX_bit_math_h_l216_c3_2748_return_output := layer0_node18_MUX_bit_math_h_l216_c3_2748_return_output;

     -- layer0_node27_MUX[bit_math_h_l315_c3_5c0f] LATENCY=0
     -- Inputs
     layer0_node27_MUX_bit_math_h_l315_c3_5c0f_cond <= VAR_layer0_node27_MUX_bit_math_h_l315_c3_5c0f_cond;
     layer0_node27_MUX_bit_math_h_l315_c3_5c0f_iftrue <= VAR_layer0_node27_MUX_bit_math_h_l315_c3_5c0f_iftrue;
     layer0_node27_MUX_bit_math_h_l315_c3_5c0f_iffalse <= VAR_layer0_node27_MUX_bit_math_h_l315_c3_5c0f_iffalse;
     -- Outputs
     VAR_layer0_node27_MUX_bit_math_h_l315_c3_5c0f_return_output := layer0_node27_MUX_bit_math_h_l315_c3_5c0f_return_output;

     -- layer0_node56_MUX[bit_math_h_l634_c3_ab19] LATENCY=0
     -- Inputs
     layer0_node56_MUX_bit_math_h_l634_c3_ab19_cond <= VAR_layer0_node56_MUX_bit_math_h_l634_c3_ab19_cond;
     layer0_node56_MUX_bit_math_h_l634_c3_ab19_iftrue <= VAR_layer0_node56_MUX_bit_math_h_l634_c3_ab19_iftrue;
     layer0_node56_MUX_bit_math_h_l634_c3_ab19_iffalse <= VAR_layer0_node56_MUX_bit_math_h_l634_c3_ab19_iffalse;
     -- Outputs
     VAR_layer0_node56_MUX_bit_math_h_l634_c3_ab19_return_output := layer0_node56_MUX_bit_math_h_l634_c3_ab19_return_output;

     -- layer0_node40_MUX[bit_math_h_l458_c3_c977] LATENCY=0
     -- Inputs
     layer0_node40_MUX_bit_math_h_l458_c3_c977_cond <= VAR_layer0_node40_MUX_bit_math_h_l458_c3_c977_cond;
     layer0_node40_MUX_bit_math_h_l458_c3_c977_iftrue <= VAR_layer0_node40_MUX_bit_math_h_l458_c3_c977_iftrue;
     layer0_node40_MUX_bit_math_h_l458_c3_c977_iffalse <= VAR_layer0_node40_MUX_bit_math_h_l458_c3_c977_iffalse;
     -- Outputs
     VAR_layer0_node40_MUX_bit_math_h_l458_c3_c977_return_output := layer0_node40_MUX_bit_math_h_l458_c3_c977_return_output;

     -- layer0_node50_MUX[bit_math_h_l568_c3_4522] LATENCY=0
     -- Inputs
     layer0_node50_MUX_bit_math_h_l568_c3_4522_cond <= VAR_layer0_node50_MUX_bit_math_h_l568_c3_4522_cond;
     layer0_node50_MUX_bit_math_h_l568_c3_4522_iftrue <= VAR_layer0_node50_MUX_bit_math_h_l568_c3_4522_iftrue;
     layer0_node50_MUX_bit_math_h_l568_c3_4522_iffalse <= VAR_layer0_node50_MUX_bit_math_h_l568_c3_4522_iffalse;
     -- Outputs
     VAR_layer0_node50_MUX_bit_math_h_l568_c3_4522_return_output := layer0_node50_MUX_bit_math_h_l568_c3_4522_return_output;

     -- layer0_node29_MUX[bit_math_h_l337_c3_cbb8] LATENCY=0
     -- Inputs
     layer0_node29_MUX_bit_math_h_l337_c3_cbb8_cond <= VAR_layer0_node29_MUX_bit_math_h_l337_c3_cbb8_cond;
     layer0_node29_MUX_bit_math_h_l337_c3_cbb8_iftrue <= VAR_layer0_node29_MUX_bit_math_h_l337_c3_cbb8_iftrue;
     layer0_node29_MUX_bit_math_h_l337_c3_cbb8_iffalse <= VAR_layer0_node29_MUX_bit_math_h_l337_c3_cbb8_iffalse;
     -- Outputs
     VAR_layer0_node29_MUX_bit_math_h_l337_c3_cbb8_return_output := layer0_node29_MUX_bit_math_h_l337_c3_cbb8_return_output;

     -- layer0_node3_MUX[bit_math_h_l51_c3_b336] LATENCY=0
     -- Inputs
     layer0_node3_MUX_bit_math_h_l51_c3_b336_cond <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_b336_cond;
     layer0_node3_MUX_bit_math_h_l51_c3_b336_iftrue <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_b336_iftrue;
     layer0_node3_MUX_bit_math_h_l51_c3_b336_iffalse <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_b336_iffalse;
     -- Outputs
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_b336_return_output := layer0_node3_MUX_bit_math_h_l51_c3_b336_return_output;

     -- layer0_node37_MUX[bit_math_h_l425_c3_2485] LATENCY=0
     -- Inputs
     layer0_node37_MUX_bit_math_h_l425_c3_2485_cond <= VAR_layer0_node37_MUX_bit_math_h_l425_c3_2485_cond;
     layer0_node37_MUX_bit_math_h_l425_c3_2485_iftrue <= VAR_layer0_node37_MUX_bit_math_h_l425_c3_2485_iftrue;
     layer0_node37_MUX_bit_math_h_l425_c3_2485_iffalse <= VAR_layer0_node37_MUX_bit_math_h_l425_c3_2485_iffalse;
     -- Outputs
     VAR_layer0_node37_MUX_bit_math_h_l425_c3_2485_return_output := layer0_node37_MUX_bit_math_h_l425_c3_2485_return_output;

     -- layer0_node32_MUX[bit_math_h_l370_c3_3d24] LATENCY=0
     -- Inputs
     layer0_node32_MUX_bit_math_h_l370_c3_3d24_cond <= VAR_layer0_node32_MUX_bit_math_h_l370_c3_3d24_cond;
     layer0_node32_MUX_bit_math_h_l370_c3_3d24_iftrue <= VAR_layer0_node32_MUX_bit_math_h_l370_c3_3d24_iftrue;
     layer0_node32_MUX_bit_math_h_l370_c3_3d24_iffalse <= VAR_layer0_node32_MUX_bit_math_h_l370_c3_3d24_iffalse;
     -- Outputs
     VAR_layer0_node32_MUX_bit_math_h_l370_c3_3d24_return_output := layer0_node32_MUX_bit_math_h_l370_c3_3d24_return_output;

     -- layer0_node53_MUX[bit_math_h_l601_c3_6dc2] LATENCY=0
     -- Inputs
     layer0_node53_MUX_bit_math_h_l601_c3_6dc2_cond <= VAR_layer0_node53_MUX_bit_math_h_l601_c3_6dc2_cond;
     layer0_node53_MUX_bit_math_h_l601_c3_6dc2_iftrue <= VAR_layer0_node53_MUX_bit_math_h_l601_c3_6dc2_iftrue;
     layer0_node53_MUX_bit_math_h_l601_c3_6dc2_iffalse <= VAR_layer0_node53_MUX_bit_math_h_l601_c3_6dc2_iffalse;
     -- Outputs
     VAR_layer0_node53_MUX_bit_math_h_l601_c3_6dc2_return_output := layer0_node53_MUX_bit_math_h_l601_c3_6dc2_return_output;

     -- layer0_node46_MUX[bit_math_h_l524_c3_4ef5] LATENCY=0
     -- Inputs
     layer0_node46_MUX_bit_math_h_l524_c3_4ef5_cond <= VAR_layer0_node46_MUX_bit_math_h_l524_c3_4ef5_cond;
     layer0_node46_MUX_bit_math_h_l524_c3_4ef5_iftrue <= VAR_layer0_node46_MUX_bit_math_h_l524_c3_4ef5_iftrue;
     layer0_node46_MUX_bit_math_h_l524_c3_4ef5_iffalse <= VAR_layer0_node46_MUX_bit_math_h_l524_c3_4ef5_iffalse;
     -- Outputs
     VAR_layer0_node46_MUX_bit_math_h_l524_c3_4ef5_return_output := layer0_node46_MUX_bit_math_h_l524_c3_4ef5_return_output;

     -- Submodule level 2
     VAR_layer1_node0_MUX_bit_math_h_l728_c3_2ff0_iffalse := VAR_layer0_node0_MUX_bit_math_h_l18_c3_5c06_return_output;
     VAR_layer1_node5_MUX_bit_math_h_l783_c3_7ab9_iffalse := VAR_layer0_node10_MUX_bit_math_h_l128_c3_0e6c_return_output;
     VAR_layer1_node5_MUX_bit_math_h_l783_c3_7ab9_iftrue := VAR_layer0_node11_MUX_bit_math_h_l139_c3_3ab9_return_output;
     VAR_layer1_node6_MUX_bit_math_h_l794_c3_1dbe_iffalse := VAR_layer0_node12_MUX_bit_math_h_l150_c3_e611_return_output;
     VAR_layer1_node6_MUX_bit_math_h_l794_c3_1dbe_iftrue := VAR_layer0_node13_MUX_bit_math_h_l161_c3_e037_return_output;
     VAR_layer1_node7_MUX_bit_math_h_l805_c3_6dfe_iffalse := VAR_layer0_node14_MUX_bit_math_h_l172_c3_ad25_return_output;
     VAR_layer1_node7_MUX_bit_math_h_l805_c3_6dfe_iftrue := VAR_layer0_node15_MUX_bit_math_h_l183_c3_dacd_return_output;
     VAR_layer1_node8_MUX_bit_math_h_l816_c3_5d19_iffalse := VAR_layer0_node16_MUX_bit_math_h_l194_c3_5393_return_output;
     VAR_layer1_node8_MUX_bit_math_h_l816_c3_5d19_iftrue := VAR_layer0_node17_MUX_bit_math_h_l205_c3_4246_return_output;
     VAR_layer1_node9_MUX_bit_math_h_l827_c3_fe3d_iffalse := VAR_layer0_node18_MUX_bit_math_h_l216_c3_2748_return_output;
     VAR_layer1_node9_MUX_bit_math_h_l827_c3_fe3d_iftrue := VAR_layer0_node19_MUX_bit_math_h_l227_c3_1dae_return_output;
     VAR_layer1_node0_MUX_bit_math_h_l728_c3_2ff0_iftrue := VAR_layer0_node1_MUX_bit_math_h_l29_c3_fa46_return_output;
     VAR_layer1_node10_MUX_bit_math_h_l838_c3_cc59_iffalse := VAR_layer0_node20_MUX_bit_math_h_l238_c3_e7c7_return_output;
     VAR_layer1_node10_MUX_bit_math_h_l838_c3_cc59_iftrue := VAR_layer0_node21_MUX_bit_math_h_l249_c3_8f8c_return_output;
     VAR_layer1_node11_MUX_bit_math_h_l849_c3_6ba8_iffalse := VAR_layer0_node22_MUX_bit_math_h_l260_c3_321e_return_output;
     VAR_layer1_node11_MUX_bit_math_h_l849_c3_6ba8_iftrue := VAR_layer0_node23_MUX_bit_math_h_l271_c3_86c3_return_output;
     VAR_layer1_node12_MUX_bit_math_h_l860_c3_e057_iffalse := VAR_layer0_node24_MUX_bit_math_h_l282_c3_2992_return_output;
     VAR_layer1_node12_MUX_bit_math_h_l860_c3_e057_iftrue := VAR_layer0_node25_MUX_bit_math_h_l293_c3_ece2_return_output;
     VAR_layer1_node13_MUX_bit_math_h_l871_c3_aad3_iffalse := VAR_layer0_node26_MUX_bit_math_h_l304_c3_7f9b_return_output;
     VAR_layer1_node13_MUX_bit_math_h_l871_c3_aad3_iftrue := VAR_layer0_node27_MUX_bit_math_h_l315_c3_5c0f_return_output;
     VAR_layer1_node14_MUX_bit_math_h_l882_c3_0d3c_iffalse := VAR_layer0_node28_MUX_bit_math_h_l326_c3_12a3_return_output;
     VAR_layer1_node14_MUX_bit_math_h_l882_c3_0d3c_iftrue := VAR_layer0_node29_MUX_bit_math_h_l337_c3_cbb8_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l739_c3_8d8d_iffalse := VAR_layer0_node2_MUX_bit_math_h_l40_c3_f68a_return_output;
     VAR_layer1_node15_MUX_bit_math_h_l893_c3_6301_iffalse := VAR_layer0_node30_MUX_bit_math_h_l348_c3_8c5c_return_output;
     VAR_layer1_node15_MUX_bit_math_h_l893_c3_6301_iftrue := VAR_layer0_node31_MUX_bit_math_h_l359_c3_d6b9_return_output;
     VAR_layer1_node16_MUX_bit_math_h_l904_c3_60f0_iffalse := VAR_layer0_node32_MUX_bit_math_h_l370_c3_3d24_return_output;
     VAR_layer1_node16_MUX_bit_math_h_l904_c3_60f0_iftrue := VAR_layer0_node33_MUX_bit_math_h_l381_c3_bdd0_return_output;
     VAR_layer1_node17_MUX_bit_math_h_l915_c3_d47f_iffalse := VAR_layer0_node34_MUX_bit_math_h_l392_c3_f617_return_output;
     VAR_layer1_node17_MUX_bit_math_h_l915_c3_d47f_iftrue := VAR_layer0_node35_MUX_bit_math_h_l403_c3_683e_return_output;
     VAR_layer1_node18_MUX_bit_math_h_l926_c3_678f_iffalse := VAR_layer0_node36_MUX_bit_math_h_l414_c3_cd2c_return_output;
     VAR_layer1_node18_MUX_bit_math_h_l926_c3_678f_iftrue := VAR_layer0_node37_MUX_bit_math_h_l425_c3_2485_return_output;
     VAR_layer1_node19_MUX_bit_math_h_l937_c3_eb8f_iffalse := VAR_layer0_node38_MUX_bit_math_h_l436_c3_c940_return_output;
     VAR_layer1_node19_MUX_bit_math_h_l937_c3_eb8f_iftrue := VAR_layer0_node39_MUX_bit_math_h_l447_c3_b150_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l739_c3_8d8d_iftrue := VAR_layer0_node3_MUX_bit_math_h_l51_c3_b336_return_output;
     VAR_layer1_node20_MUX_bit_math_h_l948_c3_588a_iffalse := VAR_layer0_node40_MUX_bit_math_h_l458_c3_c977_return_output;
     VAR_layer1_node20_MUX_bit_math_h_l948_c3_588a_iftrue := VAR_layer0_node41_MUX_bit_math_h_l469_c3_b3bf_return_output;
     VAR_layer1_node21_MUX_bit_math_h_l959_c3_1823_iffalse := VAR_layer0_node42_MUX_bit_math_h_l480_c3_c677_return_output;
     VAR_layer1_node21_MUX_bit_math_h_l959_c3_1823_iftrue := VAR_layer0_node43_MUX_bit_math_h_l491_c3_2838_return_output;
     VAR_layer1_node22_MUX_bit_math_h_l970_c3_6904_iffalse := VAR_layer0_node44_MUX_bit_math_h_l502_c3_6b96_return_output;
     VAR_layer1_node22_MUX_bit_math_h_l970_c3_6904_iftrue := VAR_layer0_node45_MUX_bit_math_h_l513_c3_b86e_return_output;
     VAR_layer1_node23_MUX_bit_math_h_l981_c3_f890_iffalse := VAR_layer0_node46_MUX_bit_math_h_l524_c3_4ef5_return_output;
     VAR_layer1_node23_MUX_bit_math_h_l981_c3_f890_iftrue := VAR_layer0_node47_MUX_bit_math_h_l535_c3_21f3_return_output;
     VAR_layer1_node24_MUX_bit_math_h_l992_c3_4e65_iffalse := VAR_layer0_node48_MUX_bit_math_h_l546_c3_5be4_return_output;
     VAR_layer1_node24_MUX_bit_math_h_l992_c3_4e65_iftrue := VAR_layer0_node49_MUX_bit_math_h_l557_c3_3410_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l750_c3_7ed6_iffalse := VAR_layer0_node4_MUX_bit_math_h_l62_c3_07e7_return_output;
     VAR_layer1_node25_MUX_bit_math_h_l1003_c3_f943_iffalse := VAR_layer0_node50_MUX_bit_math_h_l568_c3_4522_return_output;
     VAR_layer1_node25_MUX_bit_math_h_l1003_c3_f943_iftrue := VAR_layer0_node51_MUX_bit_math_h_l579_c3_8398_return_output;
     VAR_layer1_node26_MUX_bit_math_h_l1014_c3_aa20_iffalse := VAR_layer0_node52_MUX_bit_math_h_l590_c3_6d3d_return_output;
     VAR_layer1_node26_MUX_bit_math_h_l1014_c3_aa20_iftrue := VAR_layer0_node53_MUX_bit_math_h_l601_c3_6dc2_return_output;
     VAR_layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_iffalse := VAR_layer0_node54_MUX_bit_math_h_l612_c3_cab9_return_output;
     VAR_layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_iftrue := VAR_layer0_node55_MUX_bit_math_h_l623_c3_2e5e_return_output;
     VAR_layer1_node28_MUX_bit_math_h_l1036_c3_85a0_iffalse := VAR_layer0_node56_MUX_bit_math_h_l634_c3_ab19_return_output;
     VAR_layer1_node28_MUX_bit_math_h_l1036_c3_85a0_iftrue := VAR_layer0_node57_MUX_bit_math_h_l645_c3_cec5_return_output;
     VAR_layer1_node29_MUX_bit_math_h_l1047_c3_953f_iffalse := VAR_layer0_node58_MUX_bit_math_h_l656_c3_312b_return_output;
     VAR_layer1_node29_MUX_bit_math_h_l1047_c3_953f_iftrue := VAR_layer0_node59_MUX_bit_math_h_l667_c3_672d_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l750_c3_7ed6_iftrue := VAR_layer0_node5_MUX_bit_math_h_l73_c3_282b_return_output;
     VAR_layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_iffalse := VAR_layer0_node60_MUX_bit_math_h_l678_c3_9a42_return_output;
     VAR_layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_iftrue := VAR_layer0_node61_MUX_bit_math_h_l689_c3_be95_return_output;
     VAR_layer1_node31_MUX_bit_math_h_l1069_c3_82fc_iffalse := VAR_layer0_node62_MUX_bit_math_h_l700_c3_8a98_return_output;
     VAR_layer1_node31_MUX_bit_math_h_l1069_c3_82fc_iftrue := VAR_layer0_node63_MUX_bit_math_h_l711_c3_45fc_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l761_c3_68af_iffalse := VAR_layer0_node6_MUX_bit_math_h_l84_c3_62f1_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l761_c3_68af_iftrue := VAR_layer0_node7_MUX_bit_math_h_l95_c3_567b_return_output;
     VAR_layer1_node4_MUX_bit_math_h_l772_c3_e8c5_iffalse := VAR_layer0_node8_MUX_bit_math_h_l106_c3_47e5_return_output;
     VAR_layer1_node4_MUX_bit_math_h_l772_c3_e8c5_iftrue := VAR_layer0_node9_MUX_bit_math_h_l117_c3_f097_return_output;
     -- layer1_node30_MUX[bit_math_h_l1058_c3_c3ba] LATENCY=0
     -- Inputs
     layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_cond <= VAR_layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_cond;
     layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_iftrue <= VAR_layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_iftrue;
     layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_iffalse <= VAR_layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_iffalse;
     -- Outputs
     VAR_layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_return_output := layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_return_output;

     -- layer1_node7_MUX[bit_math_h_l805_c3_6dfe] LATENCY=0
     -- Inputs
     layer1_node7_MUX_bit_math_h_l805_c3_6dfe_cond <= VAR_layer1_node7_MUX_bit_math_h_l805_c3_6dfe_cond;
     layer1_node7_MUX_bit_math_h_l805_c3_6dfe_iftrue <= VAR_layer1_node7_MUX_bit_math_h_l805_c3_6dfe_iftrue;
     layer1_node7_MUX_bit_math_h_l805_c3_6dfe_iffalse <= VAR_layer1_node7_MUX_bit_math_h_l805_c3_6dfe_iffalse;
     -- Outputs
     VAR_layer1_node7_MUX_bit_math_h_l805_c3_6dfe_return_output := layer1_node7_MUX_bit_math_h_l805_c3_6dfe_return_output;

     -- layer1_node13_MUX[bit_math_h_l871_c3_aad3] LATENCY=0
     -- Inputs
     layer1_node13_MUX_bit_math_h_l871_c3_aad3_cond <= VAR_layer1_node13_MUX_bit_math_h_l871_c3_aad3_cond;
     layer1_node13_MUX_bit_math_h_l871_c3_aad3_iftrue <= VAR_layer1_node13_MUX_bit_math_h_l871_c3_aad3_iftrue;
     layer1_node13_MUX_bit_math_h_l871_c3_aad3_iffalse <= VAR_layer1_node13_MUX_bit_math_h_l871_c3_aad3_iffalse;
     -- Outputs
     VAR_layer1_node13_MUX_bit_math_h_l871_c3_aad3_return_output := layer1_node13_MUX_bit_math_h_l871_c3_aad3_return_output;

     -- layer1_node31_MUX[bit_math_h_l1069_c3_82fc] LATENCY=0
     -- Inputs
     layer1_node31_MUX_bit_math_h_l1069_c3_82fc_cond <= VAR_layer1_node31_MUX_bit_math_h_l1069_c3_82fc_cond;
     layer1_node31_MUX_bit_math_h_l1069_c3_82fc_iftrue <= VAR_layer1_node31_MUX_bit_math_h_l1069_c3_82fc_iftrue;
     layer1_node31_MUX_bit_math_h_l1069_c3_82fc_iffalse <= VAR_layer1_node31_MUX_bit_math_h_l1069_c3_82fc_iffalse;
     -- Outputs
     VAR_layer1_node31_MUX_bit_math_h_l1069_c3_82fc_return_output := layer1_node31_MUX_bit_math_h_l1069_c3_82fc_return_output;

     -- layer1_node5_MUX[bit_math_h_l783_c3_7ab9] LATENCY=0
     -- Inputs
     layer1_node5_MUX_bit_math_h_l783_c3_7ab9_cond <= VAR_layer1_node5_MUX_bit_math_h_l783_c3_7ab9_cond;
     layer1_node5_MUX_bit_math_h_l783_c3_7ab9_iftrue <= VAR_layer1_node5_MUX_bit_math_h_l783_c3_7ab9_iftrue;
     layer1_node5_MUX_bit_math_h_l783_c3_7ab9_iffalse <= VAR_layer1_node5_MUX_bit_math_h_l783_c3_7ab9_iffalse;
     -- Outputs
     VAR_layer1_node5_MUX_bit_math_h_l783_c3_7ab9_return_output := layer1_node5_MUX_bit_math_h_l783_c3_7ab9_return_output;

     -- layer1_node8_MUX[bit_math_h_l816_c3_5d19] LATENCY=0
     -- Inputs
     layer1_node8_MUX_bit_math_h_l816_c3_5d19_cond <= VAR_layer1_node8_MUX_bit_math_h_l816_c3_5d19_cond;
     layer1_node8_MUX_bit_math_h_l816_c3_5d19_iftrue <= VAR_layer1_node8_MUX_bit_math_h_l816_c3_5d19_iftrue;
     layer1_node8_MUX_bit_math_h_l816_c3_5d19_iffalse <= VAR_layer1_node8_MUX_bit_math_h_l816_c3_5d19_iffalse;
     -- Outputs
     VAR_layer1_node8_MUX_bit_math_h_l816_c3_5d19_return_output := layer1_node8_MUX_bit_math_h_l816_c3_5d19_return_output;

     -- layer1_node11_MUX[bit_math_h_l849_c3_6ba8] LATENCY=0
     -- Inputs
     layer1_node11_MUX_bit_math_h_l849_c3_6ba8_cond <= VAR_layer1_node11_MUX_bit_math_h_l849_c3_6ba8_cond;
     layer1_node11_MUX_bit_math_h_l849_c3_6ba8_iftrue <= VAR_layer1_node11_MUX_bit_math_h_l849_c3_6ba8_iftrue;
     layer1_node11_MUX_bit_math_h_l849_c3_6ba8_iffalse <= VAR_layer1_node11_MUX_bit_math_h_l849_c3_6ba8_iffalse;
     -- Outputs
     VAR_layer1_node11_MUX_bit_math_h_l849_c3_6ba8_return_output := layer1_node11_MUX_bit_math_h_l849_c3_6ba8_return_output;

     -- layer1_node17_MUX[bit_math_h_l915_c3_d47f] LATENCY=0
     -- Inputs
     layer1_node17_MUX_bit_math_h_l915_c3_d47f_cond <= VAR_layer1_node17_MUX_bit_math_h_l915_c3_d47f_cond;
     layer1_node17_MUX_bit_math_h_l915_c3_d47f_iftrue <= VAR_layer1_node17_MUX_bit_math_h_l915_c3_d47f_iftrue;
     layer1_node17_MUX_bit_math_h_l915_c3_d47f_iffalse <= VAR_layer1_node17_MUX_bit_math_h_l915_c3_d47f_iffalse;
     -- Outputs
     VAR_layer1_node17_MUX_bit_math_h_l915_c3_d47f_return_output := layer1_node17_MUX_bit_math_h_l915_c3_d47f_return_output;

     -- layer1_node19_MUX[bit_math_h_l937_c3_eb8f] LATENCY=0
     -- Inputs
     layer1_node19_MUX_bit_math_h_l937_c3_eb8f_cond <= VAR_layer1_node19_MUX_bit_math_h_l937_c3_eb8f_cond;
     layer1_node19_MUX_bit_math_h_l937_c3_eb8f_iftrue <= VAR_layer1_node19_MUX_bit_math_h_l937_c3_eb8f_iftrue;
     layer1_node19_MUX_bit_math_h_l937_c3_eb8f_iffalse <= VAR_layer1_node19_MUX_bit_math_h_l937_c3_eb8f_iffalse;
     -- Outputs
     VAR_layer1_node19_MUX_bit_math_h_l937_c3_eb8f_return_output := layer1_node19_MUX_bit_math_h_l937_c3_eb8f_return_output;

     -- layer1_node3_MUX[bit_math_h_l761_c3_68af] LATENCY=0
     -- Inputs
     layer1_node3_MUX_bit_math_h_l761_c3_68af_cond <= VAR_layer1_node3_MUX_bit_math_h_l761_c3_68af_cond;
     layer1_node3_MUX_bit_math_h_l761_c3_68af_iftrue <= VAR_layer1_node3_MUX_bit_math_h_l761_c3_68af_iftrue;
     layer1_node3_MUX_bit_math_h_l761_c3_68af_iffalse <= VAR_layer1_node3_MUX_bit_math_h_l761_c3_68af_iffalse;
     -- Outputs
     VAR_layer1_node3_MUX_bit_math_h_l761_c3_68af_return_output := layer1_node3_MUX_bit_math_h_l761_c3_68af_return_output;

     -- layer1_node14_MUX[bit_math_h_l882_c3_0d3c] LATENCY=0
     -- Inputs
     layer1_node14_MUX_bit_math_h_l882_c3_0d3c_cond <= VAR_layer1_node14_MUX_bit_math_h_l882_c3_0d3c_cond;
     layer1_node14_MUX_bit_math_h_l882_c3_0d3c_iftrue <= VAR_layer1_node14_MUX_bit_math_h_l882_c3_0d3c_iftrue;
     layer1_node14_MUX_bit_math_h_l882_c3_0d3c_iffalse <= VAR_layer1_node14_MUX_bit_math_h_l882_c3_0d3c_iffalse;
     -- Outputs
     VAR_layer1_node14_MUX_bit_math_h_l882_c3_0d3c_return_output := layer1_node14_MUX_bit_math_h_l882_c3_0d3c_return_output;

     -- layer1_node20_MUX[bit_math_h_l948_c3_588a] LATENCY=0
     -- Inputs
     layer1_node20_MUX_bit_math_h_l948_c3_588a_cond <= VAR_layer1_node20_MUX_bit_math_h_l948_c3_588a_cond;
     layer1_node20_MUX_bit_math_h_l948_c3_588a_iftrue <= VAR_layer1_node20_MUX_bit_math_h_l948_c3_588a_iftrue;
     layer1_node20_MUX_bit_math_h_l948_c3_588a_iffalse <= VAR_layer1_node20_MUX_bit_math_h_l948_c3_588a_iffalse;
     -- Outputs
     VAR_layer1_node20_MUX_bit_math_h_l948_c3_588a_return_output := layer1_node20_MUX_bit_math_h_l948_c3_588a_return_output;

     -- layer1_node15_MUX[bit_math_h_l893_c3_6301] LATENCY=0
     -- Inputs
     layer1_node15_MUX_bit_math_h_l893_c3_6301_cond <= VAR_layer1_node15_MUX_bit_math_h_l893_c3_6301_cond;
     layer1_node15_MUX_bit_math_h_l893_c3_6301_iftrue <= VAR_layer1_node15_MUX_bit_math_h_l893_c3_6301_iftrue;
     layer1_node15_MUX_bit_math_h_l893_c3_6301_iffalse <= VAR_layer1_node15_MUX_bit_math_h_l893_c3_6301_iffalse;
     -- Outputs
     VAR_layer1_node15_MUX_bit_math_h_l893_c3_6301_return_output := layer1_node15_MUX_bit_math_h_l893_c3_6301_return_output;

     -- layer1_node10_MUX[bit_math_h_l838_c3_cc59] LATENCY=0
     -- Inputs
     layer1_node10_MUX_bit_math_h_l838_c3_cc59_cond <= VAR_layer1_node10_MUX_bit_math_h_l838_c3_cc59_cond;
     layer1_node10_MUX_bit_math_h_l838_c3_cc59_iftrue <= VAR_layer1_node10_MUX_bit_math_h_l838_c3_cc59_iftrue;
     layer1_node10_MUX_bit_math_h_l838_c3_cc59_iffalse <= VAR_layer1_node10_MUX_bit_math_h_l838_c3_cc59_iffalse;
     -- Outputs
     VAR_layer1_node10_MUX_bit_math_h_l838_c3_cc59_return_output := layer1_node10_MUX_bit_math_h_l838_c3_cc59_return_output;

     -- layer1_node1_MUX[bit_math_h_l739_c3_8d8d] LATENCY=0
     -- Inputs
     layer1_node1_MUX_bit_math_h_l739_c3_8d8d_cond <= VAR_layer1_node1_MUX_bit_math_h_l739_c3_8d8d_cond;
     layer1_node1_MUX_bit_math_h_l739_c3_8d8d_iftrue <= VAR_layer1_node1_MUX_bit_math_h_l739_c3_8d8d_iftrue;
     layer1_node1_MUX_bit_math_h_l739_c3_8d8d_iffalse <= VAR_layer1_node1_MUX_bit_math_h_l739_c3_8d8d_iffalse;
     -- Outputs
     VAR_layer1_node1_MUX_bit_math_h_l739_c3_8d8d_return_output := layer1_node1_MUX_bit_math_h_l739_c3_8d8d_return_output;

     -- layer1_node9_MUX[bit_math_h_l827_c3_fe3d] LATENCY=0
     -- Inputs
     layer1_node9_MUX_bit_math_h_l827_c3_fe3d_cond <= VAR_layer1_node9_MUX_bit_math_h_l827_c3_fe3d_cond;
     layer1_node9_MUX_bit_math_h_l827_c3_fe3d_iftrue <= VAR_layer1_node9_MUX_bit_math_h_l827_c3_fe3d_iftrue;
     layer1_node9_MUX_bit_math_h_l827_c3_fe3d_iffalse <= VAR_layer1_node9_MUX_bit_math_h_l827_c3_fe3d_iffalse;
     -- Outputs
     VAR_layer1_node9_MUX_bit_math_h_l827_c3_fe3d_return_output := layer1_node9_MUX_bit_math_h_l827_c3_fe3d_return_output;

     -- layer1_node28_MUX[bit_math_h_l1036_c3_85a0] LATENCY=0
     -- Inputs
     layer1_node28_MUX_bit_math_h_l1036_c3_85a0_cond <= VAR_layer1_node28_MUX_bit_math_h_l1036_c3_85a0_cond;
     layer1_node28_MUX_bit_math_h_l1036_c3_85a0_iftrue <= VAR_layer1_node28_MUX_bit_math_h_l1036_c3_85a0_iftrue;
     layer1_node28_MUX_bit_math_h_l1036_c3_85a0_iffalse <= VAR_layer1_node28_MUX_bit_math_h_l1036_c3_85a0_iffalse;
     -- Outputs
     VAR_layer1_node28_MUX_bit_math_h_l1036_c3_85a0_return_output := layer1_node28_MUX_bit_math_h_l1036_c3_85a0_return_output;

     -- layer1_node21_MUX[bit_math_h_l959_c3_1823] LATENCY=0
     -- Inputs
     layer1_node21_MUX_bit_math_h_l959_c3_1823_cond <= VAR_layer1_node21_MUX_bit_math_h_l959_c3_1823_cond;
     layer1_node21_MUX_bit_math_h_l959_c3_1823_iftrue <= VAR_layer1_node21_MUX_bit_math_h_l959_c3_1823_iftrue;
     layer1_node21_MUX_bit_math_h_l959_c3_1823_iffalse <= VAR_layer1_node21_MUX_bit_math_h_l959_c3_1823_iffalse;
     -- Outputs
     VAR_layer1_node21_MUX_bit_math_h_l959_c3_1823_return_output := layer1_node21_MUX_bit_math_h_l959_c3_1823_return_output;

     -- layer1_node18_MUX[bit_math_h_l926_c3_678f] LATENCY=0
     -- Inputs
     layer1_node18_MUX_bit_math_h_l926_c3_678f_cond <= VAR_layer1_node18_MUX_bit_math_h_l926_c3_678f_cond;
     layer1_node18_MUX_bit_math_h_l926_c3_678f_iftrue <= VAR_layer1_node18_MUX_bit_math_h_l926_c3_678f_iftrue;
     layer1_node18_MUX_bit_math_h_l926_c3_678f_iffalse <= VAR_layer1_node18_MUX_bit_math_h_l926_c3_678f_iffalse;
     -- Outputs
     VAR_layer1_node18_MUX_bit_math_h_l926_c3_678f_return_output := layer1_node18_MUX_bit_math_h_l926_c3_678f_return_output;

     -- layer1_node16_MUX[bit_math_h_l904_c3_60f0] LATENCY=0
     -- Inputs
     layer1_node16_MUX_bit_math_h_l904_c3_60f0_cond <= VAR_layer1_node16_MUX_bit_math_h_l904_c3_60f0_cond;
     layer1_node16_MUX_bit_math_h_l904_c3_60f0_iftrue <= VAR_layer1_node16_MUX_bit_math_h_l904_c3_60f0_iftrue;
     layer1_node16_MUX_bit_math_h_l904_c3_60f0_iffalse <= VAR_layer1_node16_MUX_bit_math_h_l904_c3_60f0_iffalse;
     -- Outputs
     VAR_layer1_node16_MUX_bit_math_h_l904_c3_60f0_return_output := layer1_node16_MUX_bit_math_h_l904_c3_60f0_return_output;

     -- layer1_node2_MUX[bit_math_h_l750_c3_7ed6] LATENCY=0
     -- Inputs
     layer1_node2_MUX_bit_math_h_l750_c3_7ed6_cond <= VAR_layer1_node2_MUX_bit_math_h_l750_c3_7ed6_cond;
     layer1_node2_MUX_bit_math_h_l750_c3_7ed6_iftrue <= VAR_layer1_node2_MUX_bit_math_h_l750_c3_7ed6_iftrue;
     layer1_node2_MUX_bit_math_h_l750_c3_7ed6_iffalse <= VAR_layer1_node2_MUX_bit_math_h_l750_c3_7ed6_iffalse;
     -- Outputs
     VAR_layer1_node2_MUX_bit_math_h_l750_c3_7ed6_return_output := layer1_node2_MUX_bit_math_h_l750_c3_7ed6_return_output;

     -- layer1_node6_MUX[bit_math_h_l794_c3_1dbe] LATENCY=0
     -- Inputs
     layer1_node6_MUX_bit_math_h_l794_c3_1dbe_cond <= VAR_layer1_node6_MUX_bit_math_h_l794_c3_1dbe_cond;
     layer1_node6_MUX_bit_math_h_l794_c3_1dbe_iftrue <= VAR_layer1_node6_MUX_bit_math_h_l794_c3_1dbe_iftrue;
     layer1_node6_MUX_bit_math_h_l794_c3_1dbe_iffalse <= VAR_layer1_node6_MUX_bit_math_h_l794_c3_1dbe_iffalse;
     -- Outputs
     VAR_layer1_node6_MUX_bit_math_h_l794_c3_1dbe_return_output := layer1_node6_MUX_bit_math_h_l794_c3_1dbe_return_output;

     -- layer1_node25_MUX[bit_math_h_l1003_c3_f943] LATENCY=0
     -- Inputs
     layer1_node25_MUX_bit_math_h_l1003_c3_f943_cond <= VAR_layer1_node25_MUX_bit_math_h_l1003_c3_f943_cond;
     layer1_node25_MUX_bit_math_h_l1003_c3_f943_iftrue <= VAR_layer1_node25_MUX_bit_math_h_l1003_c3_f943_iftrue;
     layer1_node25_MUX_bit_math_h_l1003_c3_f943_iffalse <= VAR_layer1_node25_MUX_bit_math_h_l1003_c3_f943_iffalse;
     -- Outputs
     VAR_layer1_node25_MUX_bit_math_h_l1003_c3_f943_return_output := layer1_node25_MUX_bit_math_h_l1003_c3_f943_return_output;

     -- layer1_node29_MUX[bit_math_h_l1047_c3_953f] LATENCY=0
     -- Inputs
     layer1_node29_MUX_bit_math_h_l1047_c3_953f_cond <= VAR_layer1_node29_MUX_bit_math_h_l1047_c3_953f_cond;
     layer1_node29_MUX_bit_math_h_l1047_c3_953f_iftrue <= VAR_layer1_node29_MUX_bit_math_h_l1047_c3_953f_iftrue;
     layer1_node29_MUX_bit_math_h_l1047_c3_953f_iffalse <= VAR_layer1_node29_MUX_bit_math_h_l1047_c3_953f_iffalse;
     -- Outputs
     VAR_layer1_node29_MUX_bit_math_h_l1047_c3_953f_return_output := layer1_node29_MUX_bit_math_h_l1047_c3_953f_return_output;

     -- layer1_node26_MUX[bit_math_h_l1014_c3_aa20] LATENCY=0
     -- Inputs
     layer1_node26_MUX_bit_math_h_l1014_c3_aa20_cond <= VAR_layer1_node26_MUX_bit_math_h_l1014_c3_aa20_cond;
     layer1_node26_MUX_bit_math_h_l1014_c3_aa20_iftrue <= VAR_layer1_node26_MUX_bit_math_h_l1014_c3_aa20_iftrue;
     layer1_node26_MUX_bit_math_h_l1014_c3_aa20_iffalse <= VAR_layer1_node26_MUX_bit_math_h_l1014_c3_aa20_iffalse;
     -- Outputs
     VAR_layer1_node26_MUX_bit_math_h_l1014_c3_aa20_return_output := layer1_node26_MUX_bit_math_h_l1014_c3_aa20_return_output;

     -- layer1_node12_MUX[bit_math_h_l860_c3_e057] LATENCY=0
     -- Inputs
     layer1_node12_MUX_bit_math_h_l860_c3_e057_cond <= VAR_layer1_node12_MUX_bit_math_h_l860_c3_e057_cond;
     layer1_node12_MUX_bit_math_h_l860_c3_e057_iftrue <= VAR_layer1_node12_MUX_bit_math_h_l860_c3_e057_iftrue;
     layer1_node12_MUX_bit_math_h_l860_c3_e057_iffalse <= VAR_layer1_node12_MUX_bit_math_h_l860_c3_e057_iffalse;
     -- Outputs
     VAR_layer1_node12_MUX_bit_math_h_l860_c3_e057_return_output := layer1_node12_MUX_bit_math_h_l860_c3_e057_return_output;

     -- layer1_node24_MUX[bit_math_h_l992_c3_4e65] LATENCY=0
     -- Inputs
     layer1_node24_MUX_bit_math_h_l992_c3_4e65_cond <= VAR_layer1_node24_MUX_bit_math_h_l992_c3_4e65_cond;
     layer1_node24_MUX_bit_math_h_l992_c3_4e65_iftrue <= VAR_layer1_node24_MUX_bit_math_h_l992_c3_4e65_iftrue;
     layer1_node24_MUX_bit_math_h_l992_c3_4e65_iffalse <= VAR_layer1_node24_MUX_bit_math_h_l992_c3_4e65_iffalse;
     -- Outputs
     VAR_layer1_node24_MUX_bit_math_h_l992_c3_4e65_return_output := layer1_node24_MUX_bit_math_h_l992_c3_4e65_return_output;

     -- layer1_node0_MUX[bit_math_h_l728_c3_2ff0] LATENCY=0
     -- Inputs
     layer1_node0_MUX_bit_math_h_l728_c3_2ff0_cond <= VAR_layer1_node0_MUX_bit_math_h_l728_c3_2ff0_cond;
     layer1_node0_MUX_bit_math_h_l728_c3_2ff0_iftrue <= VAR_layer1_node0_MUX_bit_math_h_l728_c3_2ff0_iftrue;
     layer1_node0_MUX_bit_math_h_l728_c3_2ff0_iffalse <= VAR_layer1_node0_MUX_bit_math_h_l728_c3_2ff0_iffalse;
     -- Outputs
     VAR_layer1_node0_MUX_bit_math_h_l728_c3_2ff0_return_output := layer1_node0_MUX_bit_math_h_l728_c3_2ff0_return_output;

     -- layer1_node4_MUX[bit_math_h_l772_c3_e8c5] LATENCY=0
     -- Inputs
     layer1_node4_MUX_bit_math_h_l772_c3_e8c5_cond <= VAR_layer1_node4_MUX_bit_math_h_l772_c3_e8c5_cond;
     layer1_node4_MUX_bit_math_h_l772_c3_e8c5_iftrue <= VAR_layer1_node4_MUX_bit_math_h_l772_c3_e8c5_iftrue;
     layer1_node4_MUX_bit_math_h_l772_c3_e8c5_iffalse <= VAR_layer1_node4_MUX_bit_math_h_l772_c3_e8c5_iffalse;
     -- Outputs
     VAR_layer1_node4_MUX_bit_math_h_l772_c3_e8c5_return_output := layer1_node4_MUX_bit_math_h_l772_c3_e8c5_return_output;

     -- layer1_node23_MUX[bit_math_h_l981_c3_f890] LATENCY=0
     -- Inputs
     layer1_node23_MUX_bit_math_h_l981_c3_f890_cond <= VAR_layer1_node23_MUX_bit_math_h_l981_c3_f890_cond;
     layer1_node23_MUX_bit_math_h_l981_c3_f890_iftrue <= VAR_layer1_node23_MUX_bit_math_h_l981_c3_f890_iftrue;
     layer1_node23_MUX_bit_math_h_l981_c3_f890_iffalse <= VAR_layer1_node23_MUX_bit_math_h_l981_c3_f890_iffalse;
     -- Outputs
     VAR_layer1_node23_MUX_bit_math_h_l981_c3_f890_return_output := layer1_node23_MUX_bit_math_h_l981_c3_f890_return_output;

     -- layer1_node27_MUX[bit_math_h_l1025_c3_a3a3] LATENCY=0
     -- Inputs
     layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_cond <= VAR_layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_cond;
     layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_iftrue <= VAR_layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_iftrue;
     layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_iffalse <= VAR_layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_iffalse;
     -- Outputs
     VAR_layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_return_output := layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_return_output;

     -- layer1_node22_MUX[bit_math_h_l970_c3_6904] LATENCY=0
     -- Inputs
     layer1_node22_MUX_bit_math_h_l970_c3_6904_cond <= VAR_layer1_node22_MUX_bit_math_h_l970_c3_6904_cond;
     layer1_node22_MUX_bit_math_h_l970_c3_6904_iftrue <= VAR_layer1_node22_MUX_bit_math_h_l970_c3_6904_iftrue;
     layer1_node22_MUX_bit_math_h_l970_c3_6904_iffalse <= VAR_layer1_node22_MUX_bit_math_h_l970_c3_6904_iffalse;
     -- Outputs
     VAR_layer1_node22_MUX_bit_math_h_l970_c3_6904_return_output := layer1_node22_MUX_bit_math_h_l970_c3_6904_return_output;

     -- Submodule level 3
     VAR_layer2_node0_MUX_bit_math_h_l1086_c3_4e60_iffalse := VAR_layer1_node0_MUX_bit_math_h_l728_c3_2ff0_return_output;
     VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_iffalse := VAR_layer1_node10_MUX_bit_math_h_l838_c3_cc59_return_output;
     VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_iftrue := VAR_layer1_node11_MUX_bit_math_h_l849_c3_6ba8_return_output;
     VAR_layer2_node6_MUX_bit_math_h_l1152_c3_3828_iffalse := VAR_layer1_node12_MUX_bit_math_h_l860_c3_e057_return_output;
     VAR_layer2_node6_MUX_bit_math_h_l1152_c3_3828_iftrue := VAR_layer1_node13_MUX_bit_math_h_l871_c3_aad3_return_output;
     VAR_layer2_node7_MUX_bit_math_h_l1163_c3_f226_iffalse := VAR_layer1_node14_MUX_bit_math_h_l882_c3_0d3c_return_output;
     VAR_layer2_node7_MUX_bit_math_h_l1163_c3_f226_iftrue := VAR_layer1_node15_MUX_bit_math_h_l893_c3_6301_return_output;
     VAR_layer2_node8_MUX_bit_math_h_l1174_c3_49b7_iffalse := VAR_layer1_node16_MUX_bit_math_h_l904_c3_60f0_return_output;
     VAR_layer2_node8_MUX_bit_math_h_l1174_c3_49b7_iftrue := VAR_layer1_node17_MUX_bit_math_h_l915_c3_d47f_return_output;
     VAR_layer2_node9_MUX_bit_math_h_l1185_c3_934f_iffalse := VAR_layer1_node18_MUX_bit_math_h_l926_c3_678f_return_output;
     VAR_layer2_node9_MUX_bit_math_h_l1185_c3_934f_iftrue := VAR_layer1_node19_MUX_bit_math_h_l937_c3_eb8f_return_output;
     VAR_layer2_node0_MUX_bit_math_h_l1086_c3_4e60_iftrue := VAR_layer1_node1_MUX_bit_math_h_l739_c3_8d8d_return_output;
     VAR_layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_iffalse := VAR_layer1_node20_MUX_bit_math_h_l948_c3_588a_return_output;
     VAR_layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_iftrue := VAR_layer1_node21_MUX_bit_math_h_l959_c3_1823_return_output;
     VAR_layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_iffalse := VAR_layer1_node22_MUX_bit_math_h_l970_c3_6904_return_output;
     VAR_layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_iftrue := VAR_layer1_node23_MUX_bit_math_h_l981_c3_f890_return_output;
     VAR_layer2_node12_MUX_bit_math_h_l1218_c3_0726_iffalse := VAR_layer1_node24_MUX_bit_math_h_l992_c3_4e65_return_output;
     VAR_layer2_node12_MUX_bit_math_h_l1218_c3_0726_iftrue := VAR_layer1_node25_MUX_bit_math_h_l1003_c3_f943_return_output;
     VAR_layer2_node13_MUX_bit_math_h_l1229_c3_754d_iffalse := VAR_layer1_node26_MUX_bit_math_h_l1014_c3_aa20_return_output;
     VAR_layer2_node13_MUX_bit_math_h_l1229_c3_754d_iftrue := VAR_layer1_node27_MUX_bit_math_h_l1025_c3_a3a3_return_output;
     VAR_layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_iffalse := VAR_layer1_node28_MUX_bit_math_h_l1036_c3_85a0_return_output;
     VAR_layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_iftrue := VAR_layer1_node29_MUX_bit_math_h_l1047_c3_953f_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l1097_c3_12bb_iffalse := VAR_layer1_node2_MUX_bit_math_h_l750_c3_7ed6_return_output;
     VAR_layer2_node15_MUX_bit_math_h_l1251_c3_57b2_iffalse := VAR_layer1_node30_MUX_bit_math_h_l1058_c3_c3ba_return_output;
     VAR_layer2_node15_MUX_bit_math_h_l1251_c3_57b2_iftrue := VAR_layer1_node31_MUX_bit_math_h_l1069_c3_82fc_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l1097_c3_12bb_iftrue := VAR_layer1_node3_MUX_bit_math_h_l761_c3_68af_return_output;
     VAR_layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_iffalse := VAR_layer1_node4_MUX_bit_math_h_l772_c3_e8c5_return_output;
     VAR_layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_iftrue := VAR_layer1_node5_MUX_bit_math_h_l783_c3_7ab9_return_output;
     VAR_layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_iffalse := VAR_layer1_node6_MUX_bit_math_h_l794_c3_1dbe_return_output;
     VAR_layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_iftrue := VAR_layer1_node7_MUX_bit_math_h_l805_c3_6dfe_return_output;
     VAR_layer2_node4_MUX_bit_math_h_l1130_c3_3de0_iffalse := VAR_layer1_node8_MUX_bit_math_h_l816_c3_5d19_return_output;
     VAR_layer2_node4_MUX_bit_math_h_l1130_c3_3de0_iftrue := VAR_layer1_node9_MUX_bit_math_h_l827_c3_fe3d_return_output;
     -- layer2_node13_MUX[bit_math_h_l1229_c3_754d] LATENCY=0
     -- Inputs
     layer2_node13_MUX_bit_math_h_l1229_c3_754d_cond <= VAR_layer2_node13_MUX_bit_math_h_l1229_c3_754d_cond;
     layer2_node13_MUX_bit_math_h_l1229_c3_754d_iftrue <= VAR_layer2_node13_MUX_bit_math_h_l1229_c3_754d_iftrue;
     layer2_node13_MUX_bit_math_h_l1229_c3_754d_iffalse <= VAR_layer2_node13_MUX_bit_math_h_l1229_c3_754d_iffalse;
     -- Outputs
     VAR_layer2_node13_MUX_bit_math_h_l1229_c3_754d_return_output := layer2_node13_MUX_bit_math_h_l1229_c3_754d_return_output;

     -- layer2_node7_MUX[bit_math_h_l1163_c3_f226] LATENCY=0
     -- Inputs
     layer2_node7_MUX_bit_math_h_l1163_c3_f226_cond <= VAR_layer2_node7_MUX_bit_math_h_l1163_c3_f226_cond;
     layer2_node7_MUX_bit_math_h_l1163_c3_f226_iftrue <= VAR_layer2_node7_MUX_bit_math_h_l1163_c3_f226_iftrue;
     layer2_node7_MUX_bit_math_h_l1163_c3_f226_iffalse <= VAR_layer2_node7_MUX_bit_math_h_l1163_c3_f226_iffalse;
     -- Outputs
     VAR_layer2_node7_MUX_bit_math_h_l1163_c3_f226_return_output := layer2_node7_MUX_bit_math_h_l1163_c3_f226_return_output;

     -- layer2_node12_MUX[bit_math_h_l1218_c3_0726] LATENCY=0
     -- Inputs
     layer2_node12_MUX_bit_math_h_l1218_c3_0726_cond <= VAR_layer2_node12_MUX_bit_math_h_l1218_c3_0726_cond;
     layer2_node12_MUX_bit_math_h_l1218_c3_0726_iftrue <= VAR_layer2_node12_MUX_bit_math_h_l1218_c3_0726_iftrue;
     layer2_node12_MUX_bit_math_h_l1218_c3_0726_iffalse <= VAR_layer2_node12_MUX_bit_math_h_l1218_c3_0726_iffalse;
     -- Outputs
     VAR_layer2_node12_MUX_bit_math_h_l1218_c3_0726_return_output := layer2_node12_MUX_bit_math_h_l1218_c3_0726_return_output;

     -- layer2_node9_MUX[bit_math_h_l1185_c3_934f] LATENCY=0
     -- Inputs
     layer2_node9_MUX_bit_math_h_l1185_c3_934f_cond <= VAR_layer2_node9_MUX_bit_math_h_l1185_c3_934f_cond;
     layer2_node9_MUX_bit_math_h_l1185_c3_934f_iftrue <= VAR_layer2_node9_MUX_bit_math_h_l1185_c3_934f_iftrue;
     layer2_node9_MUX_bit_math_h_l1185_c3_934f_iffalse <= VAR_layer2_node9_MUX_bit_math_h_l1185_c3_934f_iffalse;
     -- Outputs
     VAR_layer2_node9_MUX_bit_math_h_l1185_c3_934f_return_output := layer2_node9_MUX_bit_math_h_l1185_c3_934f_return_output;

     -- layer2_node3_MUX[bit_math_h_l1119_c3_8c7b] LATENCY=0
     -- Inputs
     layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_cond <= VAR_layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_cond;
     layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_iftrue <= VAR_layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_iftrue;
     layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_iffalse <= VAR_layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_iffalse;
     -- Outputs
     VAR_layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_return_output := layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_return_output;

     -- layer2_node10_MUX[bit_math_h_l1196_c3_3f7c] LATENCY=0
     -- Inputs
     layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_cond <= VAR_layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_cond;
     layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_iftrue <= VAR_layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_iftrue;
     layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_iffalse <= VAR_layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_iffalse;
     -- Outputs
     VAR_layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_return_output := layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_return_output;

     -- layer2_node14_MUX[bit_math_h_l1240_c3_2b9a] LATENCY=0
     -- Inputs
     layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_cond <= VAR_layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_cond;
     layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_iftrue <= VAR_layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_iftrue;
     layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_iffalse <= VAR_layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_iffalse;
     -- Outputs
     VAR_layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_return_output := layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_return_output;

     -- layer2_node15_MUX[bit_math_h_l1251_c3_57b2] LATENCY=0
     -- Inputs
     layer2_node15_MUX_bit_math_h_l1251_c3_57b2_cond <= VAR_layer2_node15_MUX_bit_math_h_l1251_c3_57b2_cond;
     layer2_node15_MUX_bit_math_h_l1251_c3_57b2_iftrue <= VAR_layer2_node15_MUX_bit_math_h_l1251_c3_57b2_iftrue;
     layer2_node15_MUX_bit_math_h_l1251_c3_57b2_iffalse <= VAR_layer2_node15_MUX_bit_math_h_l1251_c3_57b2_iffalse;
     -- Outputs
     VAR_layer2_node15_MUX_bit_math_h_l1251_c3_57b2_return_output := layer2_node15_MUX_bit_math_h_l1251_c3_57b2_return_output;

     -- layer2_node8_MUX[bit_math_h_l1174_c3_49b7] LATENCY=0
     -- Inputs
     layer2_node8_MUX_bit_math_h_l1174_c3_49b7_cond <= VAR_layer2_node8_MUX_bit_math_h_l1174_c3_49b7_cond;
     layer2_node8_MUX_bit_math_h_l1174_c3_49b7_iftrue <= VAR_layer2_node8_MUX_bit_math_h_l1174_c3_49b7_iftrue;
     layer2_node8_MUX_bit_math_h_l1174_c3_49b7_iffalse <= VAR_layer2_node8_MUX_bit_math_h_l1174_c3_49b7_iffalse;
     -- Outputs
     VAR_layer2_node8_MUX_bit_math_h_l1174_c3_49b7_return_output := layer2_node8_MUX_bit_math_h_l1174_c3_49b7_return_output;

     -- layer2_node0_MUX[bit_math_h_l1086_c3_4e60] LATENCY=0
     -- Inputs
     layer2_node0_MUX_bit_math_h_l1086_c3_4e60_cond <= VAR_layer2_node0_MUX_bit_math_h_l1086_c3_4e60_cond;
     layer2_node0_MUX_bit_math_h_l1086_c3_4e60_iftrue <= VAR_layer2_node0_MUX_bit_math_h_l1086_c3_4e60_iftrue;
     layer2_node0_MUX_bit_math_h_l1086_c3_4e60_iffalse <= VAR_layer2_node0_MUX_bit_math_h_l1086_c3_4e60_iffalse;
     -- Outputs
     VAR_layer2_node0_MUX_bit_math_h_l1086_c3_4e60_return_output := layer2_node0_MUX_bit_math_h_l1086_c3_4e60_return_output;

     -- layer2_node11_MUX[bit_math_h_l1207_c3_d0a7] LATENCY=0
     -- Inputs
     layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_cond <= VAR_layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_cond;
     layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_iftrue <= VAR_layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_iftrue;
     layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_iffalse <= VAR_layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_iffalse;
     -- Outputs
     VAR_layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_return_output := layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_return_output;

     -- layer2_node2_MUX[bit_math_h_l1108_c3_fcbb] LATENCY=0
     -- Inputs
     layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_cond <= VAR_layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_cond;
     layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_iftrue <= VAR_layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_iftrue;
     layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_iffalse <= VAR_layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_iffalse;
     -- Outputs
     VAR_layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_return_output := layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_return_output;

     -- layer2_node4_MUX[bit_math_h_l1130_c3_3de0] LATENCY=0
     -- Inputs
     layer2_node4_MUX_bit_math_h_l1130_c3_3de0_cond <= VAR_layer2_node4_MUX_bit_math_h_l1130_c3_3de0_cond;
     layer2_node4_MUX_bit_math_h_l1130_c3_3de0_iftrue <= VAR_layer2_node4_MUX_bit_math_h_l1130_c3_3de0_iftrue;
     layer2_node4_MUX_bit_math_h_l1130_c3_3de0_iffalse <= VAR_layer2_node4_MUX_bit_math_h_l1130_c3_3de0_iffalse;
     -- Outputs
     VAR_layer2_node4_MUX_bit_math_h_l1130_c3_3de0_return_output := layer2_node4_MUX_bit_math_h_l1130_c3_3de0_return_output;

     -- layer2_node1_MUX[bit_math_h_l1097_c3_12bb] LATENCY=0
     -- Inputs
     layer2_node1_MUX_bit_math_h_l1097_c3_12bb_cond <= VAR_layer2_node1_MUX_bit_math_h_l1097_c3_12bb_cond;
     layer2_node1_MUX_bit_math_h_l1097_c3_12bb_iftrue <= VAR_layer2_node1_MUX_bit_math_h_l1097_c3_12bb_iftrue;
     layer2_node1_MUX_bit_math_h_l1097_c3_12bb_iffalse <= VAR_layer2_node1_MUX_bit_math_h_l1097_c3_12bb_iffalse;
     -- Outputs
     VAR_layer2_node1_MUX_bit_math_h_l1097_c3_12bb_return_output := layer2_node1_MUX_bit_math_h_l1097_c3_12bb_return_output;

     -- layer2_node5_MUX[bit_math_h_l1141_c3_a5f6] LATENCY=0
     -- Inputs
     layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_cond <= VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_cond;
     layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_iftrue <= VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_iftrue;
     layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_iffalse <= VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_iffalse;
     -- Outputs
     VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_return_output := layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_return_output;

     -- layer2_node6_MUX[bit_math_h_l1152_c3_3828] LATENCY=0
     -- Inputs
     layer2_node6_MUX_bit_math_h_l1152_c3_3828_cond <= VAR_layer2_node6_MUX_bit_math_h_l1152_c3_3828_cond;
     layer2_node6_MUX_bit_math_h_l1152_c3_3828_iftrue <= VAR_layer2_node6_MUX_bit_math_h_l1152_c3_3828_iftrue;
     layer2_node6_MUX_bit_math_h_l1152_c3_3828_iffalse <= VAR_layer2_node6_MUX_bit_math_h_l1152_c3_3828_iffalse;
     -- Outputs
     VAR_layer2_node6_MUX_bit_math_h_l1152_c3_3828_return_output := layer2_node6_MUX_bit_math_h_l1152_c3_3828_return_output;

     -- Submodule level 4
     VAR_layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_iffalse := VAR_layer2_node0_MUX_bit_math_h_l1086_c3_4e60_return_output;
     VAR_layer3_node5_MUX_bit_math_h_l1323_c3_56dd_iffalse := VAR_layer2_node10_MUX_bit_math_h_l1196_c3_3f7c_return_output;
     VAR_layer3_node5_MUX_bit_math_h_l1323_c3_56dd_iftrue := VAR_layer2_node11_MUX_bit_math_h_l1207_c3_d0a7_return_output;
     VAR_layer3_node6_MUX_bit_math_h_l1334_c3_07bd_iffalse := VAR_layer2_node12_MUX_bit_math_h_l1218_c3_0726_return_output;
     VAR_layer3_node6_MUX_bit_math_h_l1334_c3_07bd_iftrue := VAR_layer2_node13_MUX_bit_math_h_l1229_c3_754d_return_output;
     VAR_layer3_node7_MUX_bit_math_h_l1345_c3_5a50_iffalse := VAR_layer2_node14_MUX_bit_math_h_l1240_c3_2b9a_return_output;
     VAR_layer3_node7_MUX_bit_math_h_l1345_c3_5a50_iftrue := VAR_layer2_node15_MUX_bit_math_h_l1251_c3_57b2_return_output;
     VAR_layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_iftrue := VAR_layer2_node1_MUX_bit_math_h_l1097_c3_12bb_return_output;
     VAR_layer3_node1_MUX_bit_math_h_l1279_c3_73ae_iffalse := VAR_layer2_node2_MUX_bit_math_h_l1108_c3_fcbb_return_output;
     VAR_layer3_node1_MUX_bit_math_h_l1279_c3_73ae_iftrue := VAR_layer2_node3_MUX_bit_math_h_l1119_c3_8c7b_return_output;
     VAR_layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_iffalse := VAR_layer2_node4_MUX_bit_math_h_l1130_c3_3de0_return_output;
     VAR_layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_iftrue := VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a5f6_return_output;
     VAR_layer3_node3_MUX_bit_math_h_l1301_c3_827d_iffalse := VAR_layer2_node6_MUX_bit_math_h_l1152_c3_3828_return_output;
     VAR_layer3_node3_MUX_bit_math_h_l1301_c3_827d_iftrue := VAR_layer2_node7_MUX_bit_math_h_l1163_c3_f226_return_output;
     VAR_layer3_node4_MUX_bit_math_h_l1312_c3_ca04_iffalse := VAR_layer2_node8_MUX_bit_math_h_l1174_c3_49b7_return_output;
     VAR_layer3_node4_MUX_bit_math_h_l1312_c3_ca04_iftrue := VAR_layer2_node9_MUX_bit_math_h_l1185_c3_934f_return_output;
     -- layer3_node1_MUX[bit_math_h_l1279_c3_73ae] LATENCY=0
     -- Inputs
     layer3_node1_MUX_bit_math_h_l1279_c3_73ae_cond <= VAR_layer3_node1_MUX_bit_math_h_l1279_c3_73ae_cond;
     layer3_node1_MUX_bit_math_h_l1279_c3_73ae_iftrue <= VAR_layer3_node1_MUX_bit_math_h_l1279_c3_73ae_iftrue;
     layer3_node1_MUX_bit_math_h_l1279_c3_73ae_iffalse <= VAR_layer3_node1_MUX_bit_math_h_l1279_c3_73ae_iffalse;
     -- Outputs
     VAR_layer3_node1_MUX_bit_math_h_l1279_c3_73ae_return_output := layer3_node1_MUX_bit_math_h_l1279_c3_73ae_return_output;

     -- layer3_node4_MUX[bit_math_h_l1312_c3_ca04] LATENCY=0
     -- Inputs
     layer3_node4_MUX_bit_math_h_l1312_c3_ca04_cond <= VAR_layer3_node4_MUX_bit_math_h_l1312_c3_ca04_cond;
     layer3_node4_MUX_bit_math_h_l1312_c3_ca04_iftrue <= VAR_layer3_node4_MUX_bit_math_h_l1312_c3_ca04_iftrue;
     layer3_node4_MUX_bit_math_h_l1312_c3_ca04_iffalse <= VAR_layer3_node4_MUX_bit_math_h_l1312_c3_ca04_iffalse;
     -- Outputs
     VAR_layer3_node4_MUX_bit_math_h_l1312_c3_ca04_return_output := layer3_node4_MUX_bit_math_h_l1312_c3_ca04_return_output;

     -- layer3_node6_MUX[bit_math_h_l1334_c3_07bd] LATENCY=0
     -- Inputs
     layer3_node6_MUX_bit_math_h_l1334_c3_07bd_cond <= VAR_layer3_node6_MUX_bit_math_h_l1334_c3_07bd_cond;
     layer3_node6_MUX_bit_math_h_l1334_c3_07bd_iftrue <= VAR_layer3_node6_MUX_bit_math_h_l1334_c3_07bd_iftrue;
     layer3_node6_MUX_bit_math_h_l1334_c3_07bd_iffalse <= VAR_layer3_node6_MUX_bit_math_h_l1334_c3_07bd_iffalse;
     -- Outputs
     VAR_layer3_node6_MUX_bit_math_h_l1334_c3_07bd_return_output := layer3_node6_MUX_bit_math_h_l1334_c3_07bd_return_output;

     -- layer3_node2_MUX[bit_math_h_l1290_c3_d8d2] LATENCY=0
     -- Inputs
     layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_cond <= VAR_layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_cond;
     layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_iftrue <= VAR_layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_iftrue;
     layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_iffalse <= VAR_layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_iffalse;
     -- Outputs
     VAR_layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_return_output := layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_return_output;

     -- layer3_node3_MUX[bit_math_h_l1301_c3_827d] LATENCY=0
     -- Inputs
     layer3_node3_MUX_bit_math_h_l1301_c3_827d_cond <= VAR_layer3_node3_MUX_bit_math_h_l1301_c3_827d_cond;
     layer3_node3_MUX_bit_math_h_l1301_c3_827d_iftrue <= VAR_layer3_node3_MUX_bit_math_h_l1301_c3_827d_iftrue;
     layer3_node3_MUX_bit_math_h_l1301_c3_827d_iffalse <= VAR_layer3_node3_MUX_bit_math_h_l1301_c3_827d_iffalse;
     -- Outputs
     VAR_layer3_node3_MUX_bit_math_h_l1301_c3_827d_return_output := layer3_node3_MUX_bit_math_h_l1301_c3_827d_return_output;

     -- layer3_node7_MUX[bit_math_h_l1345_c3_5a50] LATENCY=0
     -- Inputs
     layer3_node7_MUX_bit_math_h_l1345_c3_5a50_cond <= VAR_layer3_node7_MUX_bit_math_h_l1345_c3_5a50_cond;
     layer3_node7_MUX_bit_math_h_l1345_c3_5a50_iftrue <= VAR_layer3_node7_MUX_bit_math_h_l1345_c3_5a50_iftrue;
     layer3_node7_MUX_bit_math_h_l1345_c3_5a50_iffalse <= VAR_layer3_node7_MUX_bit_math_h_l1345_c3_5a50_iffalse;
     -- Outputs
     VAR_layer3_node7_MUX_bit_math_h_l1345_c3_5a50_return_output := layer3_node7_MUX_bit_math_h_l1345_c3_5a50_return_output;

     -- layer3_node5_MUX[bit_math_h_l1323_c3_56dd] LATENCY=0
     -- Inputs
     layer3_node5_MUX_bit_math_h_l1323_c3_56dd_cond <= VAR_layer3_node5_MUX_bit_math_h_l1323_c3_56dd_cond;
     layer3_node5_MUX_bit_math_h_l1323_c3_56dd_iftrue <= VAR_layer3_node5_MUX_bit_math_h_l1323_c3_56dd_iftrue;
     layer3_node5_MUX_bit_math_h_l1323_c3_56dd_iffalse <= VAR_layer3_node5_MUX_bit_math_h_l1323_c3_56dd_iffalse;
     -- Outputs
     VAR_layer3_node5_MUX_bit_math_h_l1323_c3_56dd_return_output := layer3_node5_MUX_bit_math_h_l1323_c3_56dd_return_output;

     -- layer3_node0_MUX[bit_math_h_l1268_c3_e5cc] LATENCY=0
     -- Inputs
     layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_cond <= VAR_layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_cond;
     layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_iftrue <= VAR_layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_iftrue;
     layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_iffalse <= VAR_layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_iffalse;
     -- Outputs
     VAR_layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_return_output := layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_return_output;

     -- Submodule level 5
     VAR_layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_iffalse := VAR_layer3_node0_MUX_bit_math_h_l1268_c3_e5cc_return_output;
     VAR_layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_iftrue := VAR_layer3_node1_MUX_bit_math_h_l1279_c3_73ae_return_output;
     VAR_layer4_node1_MUX_bit_math_h_l1373_c3_402b_iffalse := VAR_layer3_node2_MUX_bit_math_h_l1290_c3_d8d2_return_output;
     VAR_layer4_node1_MUX_bit_math_h_l1373_c3_402b_iftrue := VAR_layer3_node3_MUX_bit_math_h_l1301_c3_827d_return_output;
     VAR_layer4_node2_MUX_bit_math_h_l1384_c3_5f80_iffalse := VAR_layer3_node4_MUX_bit_math_h_l1312_c3_ca04_return_output;
     VAR_layer4_node2_MUX_bit_math_h_l1384_c3_5f80_iftrue := VAR_layer3_node5_MUX_bit_math_h_l1323_c3_56dd_return_output;
     VAR_layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_iffalse := VAR_layer3_node6_MUX_bit_math_h_l1334_c3_07bd_return_output;
     VAR_layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_iftrue := VAR_layer3_node7_MUX_bit_math_h_l1345_c3_5a50_return_output;
     -- layer4_node3_MUX[bit_math_h_l1395_c3_4d9c] LATENCY=0
     -- Inputs
     layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_cond <= VAR_layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_cond;
     layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_iftrue <= VAR_layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_iftrue;
     layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_iffalse <= VAR_layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_iffalse;
     -- Outputs
     VAR_layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_return_output := layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_return_output;

     -- layer4_node1_MUX[bit_math_h_l1373_c3_402b] LATENCY=0
     -- Inputs
     layer4_node1_MUX_bit_math_h_l1373_c3_402b_cond <= VAR_layer4_node1_MUX_bit_math_h_l1373_c3_402b_cond;
     layer4_node1_MUX_bit_math_h_l1373_c3_402b_iftrue <= VAR_layer4_node1_MUX_bit_math_h_l1373_c3_402b_iftrue;
     layer4_node1_MUX_bit_math_h_l1373_c3_402b_iffalse <= VAR_layer4_node1_MUX_bit_math_h_l1373_c3_402b_iffalse;
     -- Outputs
     VAR_layer4_node1_MUX_bit_math_h_l1373_c3_402b_return_output := layer4_node1_MUX_bit_math_h_l1373_c3_402b_return_output;

     -- layer4_node2_MUX[bit_math_h_l1384_c3_5f80] LATENCY=0
     -- Inputs
     layer4_node2_MUX_bit_math_h_l1384_c3_5f80_cond <= VAR_layer4_node2_MUX_bit_math_h_l1384_c3_5f80_cond;
     layer4_node2_MUX_bit_math_h_l1384_c3_5f80_iftrue <= VAR_layer4_node2_MUX_bit_math_h_l1384_c3_5f80_iftrue;
     layer4_node2_MUX_bit_math_h_l1384_c3_5f80_iffalse <= VAR_layer4_node2_MUX_bit_math_h_l1384_c3_5f80_iffalse;
     -- Outputs
     VAR_layer4_node2_MUX_bit_math_h_l1384_c3_5f80_return_output := layer4_node2_MUX_bit_math_h_l1384_c3_5f80_return_output;

     -- layer4_node0_MUX[bit_math_h_l1362_c3_f5a3] LATENCY=0
     -- Inputs
     layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_cond <= VAR_layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_cond;
     layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_iftrue <= VAR_layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_iftrue;
     layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_iffalse <= VAR_layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_iffalse;
     -- Outputs
     VAR_layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_return_output := layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_return_output;

     -- Submodule level 6
     VAR_layer5_node0_MUX_bit_math_h_l1412_c3_19e3_iffalse := VAR_layer4_node0_MUX_bit_math_h_l1362_c3_f5a3_return_output;
     VAR_layer5_node0_MUX_bit_math_h_l1412_c3_19e3_iftrue := VAR_layer4_node1_MUX_bit_math_h_l1373_c3_402b_return_output;
     VAR_layer5_node1_MUX_bit_math_h_l1423_c3_11f1_iffalse := VAR_layer4_node2_MUX_bit_math_h_l1384_c3_5f80_return_output;
     VAR_layer5_node1_MUX_bit_math_h_l1423_c3_11f1_iftrue := VAR_layer4_node3_MUX_bit_math_h_l1395_c3_4d9c_return_output;
     -- layer5_node0_MUX[bit_math_h_l1412_c3_19e3] LATENCY=0
     -- Inputs
     layer5_node0_MUX_bit_math_h_l1412_c3_19e3_cond <= VAR_layer5_node0_MUX_bit_math_h_l1412_c3_19e3_cond;
     layer5_node0_MUX_bit_math_h_l1412_c3_19e3_iftrue <= VAR_layer5_node0_MUX_bit_math_h_l1412_c3_19e3_iftrue;
     layer5_node0_MUX_bit_math_h_l1412_c3_19e3_iffalse <= VAR_layer5_node0_MUX_bit_math_h_l1412_c3_19e3_iffalse;
     -- Outputs
     VAR_layer5_node0_MUX_bit_math_h_l1412_c3_19e3_return_output := layer5_node0_MUX_bit_math_h_l1412_c3_19e3_return_output;

     -- layer5_node1_MUX[bit_math_h_l1423_c3_11f1] LATENCY=0
     -- Inputs
     layer5_node1_MUX_bit_math_h_l1423_c3_11f1_cond <= VAR_layer5_node1_MUX_bit_math_h_l1423_c3_11f1_cond;
     layer5_node1_MUX_bit_math_h_l1423_c3_11f1_iftrue <= VAR_layer5_node1_MUX_bit_math_h_l1423_c3_11f1_iftrue;
     layer5_node1_MUX_bit_math_h_l1423_c3_11f1_iffalse <= VAR_layer5_node1_MUX_bit_math_h_l1423_c3_11f1_iffalse;
     -- Outputs
     VAR_layer5_node1_MUX_bit_math_h_l1423_c3_11f1_return_output := layer5_node1_MUX_bit_math_h_l1423_c3_11f1_return_output;

     -- Submodule level 7
     VAR_layer6_node0_MUX_bit_math_h_l1440_c3_f906_iffalse := VAR_layer5_node0_MUX_bit_math_h_l1412_c3_19e3_return_output;
     VAR_layer6_node0_MUX_bit_math_h_l1440_c3_f906_iftrue := VAR_layer5_node1_MUX_bit_math_h_l1423_c3_11f1_return_output;
     -- layer6_node0_MUX[bit_math_h_l1440_c3_f906] LATENCY=0
     -- Inputs
     layer6_node0_MUX_bit_math_h_l1440_c3_f906_cond <= VAR_layer6_node0_MUX_bit_math_h_l1440_c3_f906_cond;
     layer6_node0_MUX_bit_math_h_l1440_c3_f906_iftrue <= VAR_layer6_node0_MUX_bit_math_h_l1440_c3_f906_iftrue;
     layer6_node0_MUX_bit_math_h_l1440_c3_f906_iffalse <= VAR_layer6_node0_MUX_bit_math_h_l1440_c3_f906_iffalse;
     -- Outputs
     VAR_layer6_node0_MUX_bit_math_h_l1440_c3_f906_return_output := layer6_node0_MUX_bit_math_h_l1440_c3_f906_return_output;

     -- Submodule level 8
     VAR_return_output := VAR_layer6_node0_MUX_bit_math_h_l1440_c3_f906_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
