-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity gth_0CLK_441a128d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end gth_0CLK_441a128d;
architecture arch of gth_0CLK_441a128d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1809_c6_427e]
signal BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1809_c2_ad01]
signal t8_MUX_uxn_opcodes_h_l1809_c2_ad01_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1809_c2_ad01]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1809_c2_ad01]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1809_c2_ad01]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1809_c2_ad01]
signal result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1809_c2_ad01]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1809_c2_ad01]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1809_c2_ad01]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1809_c2_ad01]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1809_c2_ad01]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output : unsigned(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l1809_c2_ad01]
signal n8_MUX_uxn_opcodes_h_l1809_c2_ad01_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1822_c11_941a]
signal BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1822_c7_ba42]
signal t8_MUX_uxn_opcodes_h_l1822_c7_ba42_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1822_c7_ba42]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1822_c7_ba42]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1822_c7_ba42]
signal result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1822_c7_ba42]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1822_c7_ba42]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output : unsigned(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l1822_c7_ba42]
signal n8_MUX_uxn_opcodes_h_l1822_c7_ba42_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1825_c11_6b04]
signal BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1825_c7_bba7]
signal t8_MUX_uxn_opcodes_h_l1825_c7_bba7_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1825_c7_bba7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1825_c7_bba7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1825_c7_bba7]
signal result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1825_c7_bba7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1825_c7_bba7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output : unsigned(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l1825_c7_bba7]
signal n8_MUX_uxn_opcodes_h_l1825_c7_bba7_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1828_c11_b4b4]
signal BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1828_c7_f8f1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1828_c7_f8f1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1828_c7_f8f1]
signal result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1828_c7_f8f1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1828_c7_f8f1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output : unsigned(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l1828_c7_f8f1]
signal n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1830_c30_20ca]
signal sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_return_output : signed(3 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1833_c21_6652]
signal BIN_OP_GT_uxn_opcodes_h_l1833_c21_6652_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1833_c21_6652_right : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1833_c21_6652_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1833_c21_1bbe]
signal MUX_uxn_opcodes_h_l1833_c21_1bbe_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1833_c21_1bbe_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1833_c21_1bbe_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1833_c21_1bbe_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_71f0( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_index_flipped := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.stack_address_sp_offset := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e
BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_left,
BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_right,
BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_return_output);

-- t8_MUX_uxn_opcodes_h_l1809_c2_ad01
t8_MUX_uxn_opcodes_h_l1809_c2_ad01 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1809_c2_ad01_cond,
t8_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue,
t8_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse,
t8_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01
result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01
result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01
result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_cond,
result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01
result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01
result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01
result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01
result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output);

-- n8_MUX_uxn_opcodes_h_l1809_c2_ad01
n8_MUX_uxn_opcodes_h_l1809_c2_ad01 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1809_c2_ad01_cond,
n8_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue,
n8_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse,
n8_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a
BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_left,
BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_right,
BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_return_output);

-- t8_MUX_uxn_opcodes_h_l1822_c7_ba42
t8_MUX_uxn_opcodes_h_l1822_c7_ba42 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1822_c7_ba42_cond,
t8_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue,
t8_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse,
t8_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42
result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42
result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42
result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_cond,
result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42
result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output);

-- n8_MUX_uxn_opcodes_h_l1822_c7_ba42
n8_MUX_uxn_opcodes_h_l1822_c7_ba42 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1822_c7_ba42_cond,
n8_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue,
n8_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse,
n8_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04
BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_left,
BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_right,
BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_return_output);

-- t8_MUX_uxn_opcodes_h_l1825_c7_bba7
t8_MUX_uxn_opcodes_h_l1825_c7_bba7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1825_c7_bba7_cond,
t8_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue,
t8_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse,
t8_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7
result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7
result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7
result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_cond,
result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7
result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output);

-- n8_MUX_uxn_opcodes_h_l1825_c7_bba7
n8_MUX_uxn_opcodes_h_l1825_c7_bba7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1825_c7_bba7_cond,
n8_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue,
n8_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse,
n8_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4
BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4_left,
BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4_right,
BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1
result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1
result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1
result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond,
result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1
result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output);

-- n8_MUX_uxn_opcodes_h_l1828_c7_f8f1
n8_MUX_uxn_opcodes_h_l1828_c7_f8f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond,
n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue,
n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse,
n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca
sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_ins,
sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_x,
sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_y,
sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1833_c21_6652
BIN_OP_GT_uxn_opcodes_h_l1833_c21_6652 : entity work.BIN_OP_GT_uint8_t_uint8_t_0CLK_380ecc95 port map (
BIN_OP_GT_uxn_opcodes_h_l1833_c21_6652_left,
BIN_OP_GT_uxn_opcodes_h_l1833_c21_6652_right,
BIN_OP_GT_uxn_opcodes_h_l1833_c21_6652_return_output);

-- MUX_uxn_opcodes_h_l1833_c21_1bbe
MUX_uxn_opcodes_h_l1833_c21_1bbe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1833_c21_1bbe_cond,
MUX_uxn_opcodes_h_l1833_c21_1bbe_iftrue,
MUX_uxn_opcodes_h_l1833_c21_1bbe_iffalse,
MUX_uxn_opcodes_h_l1833_c21_1bbe_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_return_output,
 t8_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output,
 n8_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_return_output,
 t8_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output,
 n8_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_return_output,
 t8_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output,
 n8_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output,
 n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output,
 sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1833_c21_6652_return_output,
 MUX_uxn_opcodes_h_l1833_c21_1bbe_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1809_c2_ad01_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1809_c2_ad01_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1809_c2_ad01_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1814_c3_4988 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1809_c2_ad01_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1809_c2_ad01_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1819_c3_bbf4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1809_c2_ad01_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1822_c7_ba42_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1823_c3_a31e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1822_c7_ba42_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1825_c7_bba7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1825_c7_bba7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1832_c3_7830 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1833_c21_1bbe_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_6652_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_6652_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_6652_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1833_c21_1bbe_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1833_c21_1bbe_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1833_c21_1bbe_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1825_l1809_l1828_l1822_DUPLICATE_8736_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_3ee0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_61c3_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_9641_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1825_l1828_DUPLICATE_23d7_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l1837_l1805_DUPLICATE_a345_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1832_c3_7830 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1832_c3_7830;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1833_c21_1bbe_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1833_c21_1bbe_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1823_c3_a31e := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1823_c3_a31e;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4_right := to_unsigned(3, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1814_c3_4988 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1814_c3_4988;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1819_c3_bbf4 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1819_c3_bbf4;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4_left := VAR_phase;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_6652_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_6652_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse := t8;
     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1809_c2_ad01] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1809_c2_ad01_return_output := result.is_pc_updated;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1809_c2_ad01] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1809_c2_ad01_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l1809_c6_427e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_9641 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_9641_return_output := result.is_opc_done;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1809_c2_ad01] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1809_c2_ad01_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1828_c11_b4b4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4_left;
     BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4_return_output := BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1830_c30_20ca] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_ins;
     sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_x;
     sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_return_output := sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1825_l1809_l1828_l1822_DUPLICATE_8736 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1825_l1809_l1828_l1822_DUPLICATE_8736_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1825_c11_6b04] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_left;
     BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_return_output := BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_61c3 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_61c3_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1825_l1828_DUPLICATE_23d7 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1825_l1828_DUPLICATE_23d7_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_3ee0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_3ee0_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1822_c11_941a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l1833_c21_6652] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1833_c21_6652_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_6652_left;
     BIN_OP_GT_uxn_opcodes_h_l1833_c21_6652_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_6652_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_6652_return_output := BIN_OP_GT_uxn_opcodes_h_l1833_c21_6652_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1809_c2_ad01] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1809_c2_ad01_return_output := result.is_vram_write;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1809_c2_ad01_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1809_c2_ad01_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1809_c6_427e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1822_c7_ba42_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1822_c7_ba42_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1822_c11_941a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1825_c7_bba7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1825_c7_bba7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1825_c11_6b04_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1828_c11_b4b4_return_output;
     VAR_MUX_uxn_opcodes_h_l1833_c21_1bbe_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1833_c21_6652_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_61c3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_61c3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_61c3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_9641_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_9641_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_9641_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_3ee0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_3ee0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1825_l1828_l1822_DUPLICATE_3ee0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1825_l1828_DUPLICATE_23d7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1825_l1828_DUPLICATE_23d7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1825_l1809_l1828_l1822_DUPLICATE_8736_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1825_l1809_l1828_l1822_DUPLICATE_8736_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1825_l1809_l1828_l1822_DUPLICATE_8736_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1825_l1809_l1828_l1822_DUPLICATE_8736_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1809_c2_ad01_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1809_c2_ad01_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1809_c2_ad01_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1809_c2_ad01_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1830_c30_20ca_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1828_c7_f8f1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1809_c2_ad01] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1809_c2_ad01] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output;

     -- n8_MUX[uxn_opcodes_h_l1828_c7_f8f1] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond <= VAR_n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond;
     n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue;
     n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output := n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1828_c7_f8f1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output;

     -- t8_MUX[uxn_opcodes_h_l1825_c7_bba7] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1825_c7_bba7_cond <= VAR_t8_MUX_uxn_opcodes_h_l1825_c7_bba7_cond;
     t8_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue;
     t8_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output := t8_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1828_c7_f8f1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1809_c2_ad01] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1809_c2_ad01] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1828_c7_f8f1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output;

     -- MUX[uxn_opcodes_h_l1833_c21_1bbe] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1833_c21_1bbe_cond <= VAR_MUX_uxn_opcodes_h_l1833_c21_1bbe_cond;
     MUX_uxn_opcodes_h_l1833_c21_1bbe_iftrue <= VAR_MUX_uxn_opcodes_h_l1833_c21_1bbe_iftrue;
     MUX_uxn_opcodes_h_l1833_c21_1bbe_iffalse <= VAR_MUX_uxn_opcodes_h_l1833_c21_1bbe_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1833_c21_1bbe_return_output := MUX_uxn_opcodes_h_l1833_c21_1bbe_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue := VAR_MUX_uxn_opcodes_h_l1833_c21_1bbe_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output;
     -- n8_MUX[uxn_opcodes_h_l1825_c7_bba7] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1825_c7_bba7_cond <= VAR_n8_MUX_uxn_opcodes_h_l1825_c7_bba7_cond;
     n8_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue;
     n8_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output := n8_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1825_c7_bba7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1825_c7_bba7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1825_c7_bba7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output;

     -- t8_MUX[uxn_opcodes_h_l1822_c7_ba42] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1822_c7_ba42_cond <= VAR_t8_MUX_uxn_opcodes_h_l1822_c7_ba42_cond;
     t8_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue;
     t8_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output := t8_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1825_c7_bba7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1828_c7_f8f1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output := result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1828_c7_f8f1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output;
     -- t8_MUX[uxn_opcodes_h_l1809_c2_ad01] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1809_c2_ad01_cond <= VAR_t8_MUX_uxn_opcodes_h_l1809_c2_ad01_cond;
     t8_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue;
     t8_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output := t8_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1822_c7_ba42] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1822_c7_ba42] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1822_c7_ba42] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1822_c7_ba42] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1825_c7_bba7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output := result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output;

     -- n8_MUX[uxn_opcodes_h_l1822_c7_ba42] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1822_c7_ba42_cond <= VAR_n8_MUX_uxn_opcodes_h_l1822_c7_ba42_cond;
     n8_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue;
     n8_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output := n8_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1825_c7_bba7_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1809_c2_ad01] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1809_c2_ad01] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1809_c2_ad01] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1809_c2_ad01] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1822_c7_ba42] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output := result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output;

     -- n8_MUX[uxn_opcodes_h_l1809_c2_ad01] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1809_c2_ad01_cond <= VAR_n8_MUX_uxn_opcodes_h_l1809_c2_ad01_cond;
     n8_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue;
     n8_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output := n8_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1822_c7_ba42_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1809_c2_ad01] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output := result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l1837_l1805_DUPLICATE_a345 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l1837_l1805_DUPLICATE_a345_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_71f0(
     result,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1809_c2_ad01_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l1837_l1805_DUPLICATE_a345_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l1837_l1805_DUPLICATE_a345_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
