-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 47
entity deo_0CLK_aac5017e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_device_ram_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end deo_0CLK_aac5017e;
architecture arch of deo_0CLK_aac5017e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal device_out_result : device_out_result_t := device_out_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;
signal REG_COMB_device_out_result : device_out_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l502_c6_d85c]
signal BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l509_c7_95b1]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : unsigned(0 downto 0);

-- device_out_result_MUX[uxn_opcodes_h_l502_c2_1228]
signal device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_cond : unsigned(0 downto 0);
signal device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_iftrue : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_iffalse : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_return_output : device_out_result_t;

-- n8_MUX[uxn_opcodes_h_l502_c2_1228]
signal n8_MUX_uxn_opcodes_h_l502_c2_1228_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l502_c2_1228_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l502_c2_1228_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l502_c2_1228_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l502_c2_1228]
signal result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_return_output : unsigned(7 downto 0);

-- result_vram_write_layer_MUX[uxn_opcodes_h_l502_c2_1228]
signal result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_cond : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_iftrue : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_iffalse : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l502_c2_1228]
signal result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l502_c2_1228]
signal result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_return_output : unsigned(15 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l502_c2_1228]
signal result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l502_c2_1228]
signal result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_return_output : unsigned(0 downto 0);

-- result_is_device_ram_write_MUX[uxn_opcodes_h_l502_c2_1228]
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_cond : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l502_c2_1228]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l502_c2_1228]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l502_c2_1228]
signal t8_MUX_uxn_opcodes_h_l502_c2_1228_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l502_c2_1228_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l502_c2_1228_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l502_c2_1228_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l509_c11_500d]
signal BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l512_c7_21e6]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_return_output : unsigned(0 downto 0);

-- device_out_result_MUX[uxn_opcodes_h_l509_c7_95b1]
signal device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
signal device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : device_out_result_t;

-- n8_MUX[uxn_opcodes_h_l509_c7_95b1]
signal n8_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l509_c7_95b1]
signal result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : unsigned(7 downto 0);

-- result_vram_write_layer_MUX[uxn_opcodes_h_l509_c7_95b1]
signal result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l509_c7_95b1]
signal result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l509_c7_95b1]
signal result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : unsigned(15 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l509_c7_95b1]
signal result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l509_c7_95b1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : unsigned(0 downto 0);

-- result_is_device_ram_write_MUX[uxn_opcodes_h_l509_c7_95b1]
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l509_c7_95b1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l509_c7_95b1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l509_c7_95b1]
signal t8_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l512_c11_3193]
signal BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l517_c1_4eeb]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_return_output : unsigned(0 downto 0);

-- device_out_result_MUX[uxn_opcodes_h_l512_c7_21e6]
signal device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_cond : unsigned(0 downto 0);
signal device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse : device_out_result_t;
signal device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_return_output : device_out_result_t;

-- n8_MUX[uxn_opcodes_h_l512_c7_21e6]
signal n8_MUX_uxn_opcodes_h_l512_c7_21e6_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l512_c7_21e6_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l512_c7_21e6]
signal result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_return_output : unsigned(7 downto 0);

-- result_vram_write_layer_MUX[uxn_opcodes_h_l512_c7_21e6]
signal result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_cond : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse : unsigned(0 downto 0);
signal result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l512_c7_21e6]
signal result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l512_c7_21e6]
signal result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_return_output : unsigned(15 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l512_c7_21e6]
signal result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l512_c7_21e6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_return_output : unsigned(0 downto 0);

-- result_is_device_ram_write_MUX[uxn_opcodes_h_l512_c7_21e6]
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_cond : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l512_c7_21e6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l512_c7_21e6]
signal t8_MUX_uxn_opcodes_h_l512_c7_21e6_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l512_c7_21e6_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l515_c30_e5ba]
signal sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l519_c9_614a]
signal BIN_OP_EQ_uxn_opcodes_h_l519_c9_614a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l519_c9_614a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l519_c9_614a_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l519_c9_1c10]
signal MUX_uxn_opcodes_h_l519_c9_1c10_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l519_c9_1c10_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l519_c9_1c10_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l519_c9_1c10_return_output : unsigned(7 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_h_l520_c42_ad6a]
signal BIN_OP_MINUS_uxn_opcodes_h_l520_c42_ad6a_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l520_c42_ad6a_right : unsigned(1 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l520_c42_ad6a_return_output : unsigned(7 downto 0);

-- device_out[uxn_opcodes_h_l520_c23_fa5d]
signal device_out_uxn_opcodes_h_l520_c23_fa5d_CLOCK_ENABLE : unsigned(0 downto 0);
signal device_out_uxn_opcodes_h_l520_c23_fa5d_device_address : unsigned(7 downto 0);
signal device_out_uxn_opcodes_h_l520_c23_fa5d_value : unsigned(7 downto 0);
signal device_out_uxn_opcodes_h_l520_c23_fa5d_phase : unsigned(7 downto 0);
signal device_out_uxn_opcodes_h_l520_c23_fa5d_previous_device_ram_read : unsigned(7 downto 0);
signal device_out_uxn_opcodes_h_l520_c23_fa5d_previous_ram_read : unsigned(7 downto 0);
signal device_out_uxn_opcodes_h_l520_c23_fa5d_return_output : device_out_result_t;

function CONST_REF_RD_opcode_result_t_opcode_result_t_23b1( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.vram_write_layer := ref_toks_2;
      base.is_vram_write := ref_toks_3;
      base.u16_value := ref_toks_4;
      base.device_ram_address := ref_toks_5;
      base.is_opc_done := ref_toks_6;
      base.is_device_ram_write := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.sp_relative_shift := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c
BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_left,
BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_right,
BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_return_output);

-- device_out_result_MUX_uxn_opcodes_h_l502_c2_1228
device_out_result_MUX_uxn_opcodes_h_l502_c2_1228 : entity work.MUX_uint1_t_device_out_result_t_device_out_result_t_0CLK_de264c78 port map (
device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_cond,
device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_iftrue,
device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_iffalse,
device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_return_output);

-- n8_MUX_uxn_opcodes_h_l502_c2_1228
n8_MUX_uxn_opcodes_h_l502_c2_1228 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l502_c2_1228_cond,
n8_MUX_uxn_opcodes_h_l502_c2_1228_iftrue,
n8_MUX_uxn_opcodes_h_l502_c2_1228_iffalse,
n8_MUX_uxn_opcodes_h_l502_c2_1228_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228
result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_cond,
result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_return_output);

-- result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228
result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_cond,
result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_iftrue,
result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_iffalse,
result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228
result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228
result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_cond,
result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228
result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228
result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_return_output);

-- result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228
result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_cond,
result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_iftrue,
result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_iffalse,
result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228
result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_return_output);

-- t8_MUX_uxn_opcodes_h_l502_c2_1228
t8_MUX_uxn_opcodes_h_l502_c2_1228 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l502_c2_1228_cond,
t8_MUX_uxn_opcodes_h_l502_c2_1228_iftrue,
t8_MUX_uxn_opcodes_h_l502_c2_1228_iffalse,
t8_MUX_uxn_opcodes_h_l502_c2_1228_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d
BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_left,
BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_right,
BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_return_output);

-- device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1
device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1 : entity work.MUX_uint1_t_device_out_result_t_device_out_result_t_0CLK_de264c78 port map (
device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_cond,
device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue,
device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse,
device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_return_output);

-- n8_MUX_uxn_opcodes_h_l509_c7_95b1
n8_MUX_uxn_opcodes_h_l509_c7_95b1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l509_c7_95b1_cond,
n8_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue,
n8_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse,
n8_MUX_uxn_opcodes_h_l509_c7_95b1_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1
result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_cond,
result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_return_output);

-- result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1
result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_cond,
result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue,
result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse,
result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1
result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1
result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_cond,
result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1
result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1
result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_return_output);

-- result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1
result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_cond,
result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue,
result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse,
result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1
result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_return_output);

-- t8_MUX_uxn_opcodes_h_l509_c7_95b1
t8_MUX_uxn_opcodes_h_l509_c7_95b1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l509_c7_95b1_cond,
t8_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue,
t8_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse,
t8_MUX_uxn_opcodes_h_l509_c7_95b1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193
BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_left,
BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_right,
BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_return_output);

-- device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6
device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6 : entity work.MUX_uint1_t_device_out_result_t_device_out_result_t_0CLK_de264c78 port map (
device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_cond,
device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue,
device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse,
device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_return_output);

-- n8_MUX_uxn_opcodes_h_l512_c7_21e6
n8_MUX_uxn_opcodes_h_l512_c7_21e6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l512_c7_21e6_cond,
n8_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue,
n8_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse,
n8_MUX_uxn_opcodes_h_l512_c7_21e6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6
result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_cond,
result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_return_output);

-- result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6
result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_cond,
result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue,
result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse,
result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6
result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6
result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_cond,
result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6
result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6
result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_return_output);

-- result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6
result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_cond,
result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue,
result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse,
result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6
result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_return_output);

-- t8_MUX_uxn_opcodes_h_l512_c7_21e6
t8_MUX_uxn_opcodes_h_l512_c7_21e6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l512_c7_21e6_cond,
t8_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue,
t8_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse,
t8_MUX_uxn_opcodes_h_l512_c7_21e6_return_output);

-- sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba
sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_ins,
sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_x,
sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_y,
sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l519_c9_614a
BIN_OP_EQ_uxn_opcodes_h_l519_c9_614a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l519_c9_614a_left,
BIN_OP_EQ_uxn_opcodes_h_l519_c9_614a_right,
BIN_OP_EQ_uxn_opcodes_h_l519_c9_614a_return_output);

-- MUX_uxn_opcodes_h_l519_c9_1c10
MUX_uxn_opcodes_h_l519_c9_1c10 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l519_c9_1c10_cond,
MUX_uxn_opcodes_h_l519_c9_1c10_iftrue,
MUX_uxn_opcodes_h_l519_c9_1c10_iffalse,
MUX_uxn_opcodes_h_l519_c9_1c10_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l520_c42_ad6a
BIN_OP_MINUS_uxn_opcodes_h_l520_c42_ad6a : entity work.BIN_OP_MINUS_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l520_c42_ad6a_left,
BIN_OP_MINUS_uxn_opcodes_h_l520_c42_ad6a_right,
BIN_OP_MINUS_uxn_opcodes_h_l520_c42_ad6a_return_output);

-- device_out_uxn_opcodes_h_l520_c23_fa5d
device_out_uxn_opcodes_h_l520_c23_fa5d : entity work.device_out_0CLK_95124a2a port map (
clk,
device_out_uxn_opcodes_h_l520_c23_fa5d_CLOCK_ENABLE,
device_out_uxn_opcodes_h_l520_c23_fa5d_device_address,
device_out_uxn_opcodes_h_l520_c23_fa5d_value,
device_out_uxn_opcodes_h_l520_c23_fa5d_phase,
device_out_uxn_opcodes_h_l520_c23_fa5d_previous_device_ram_read,
device_out_uxn_opcodes_h_l520_c23_fa5d_previous_ram_read,
device_out_uxn_opcodes_h_l520_c23_fa5d_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_device_ram_read,
 previous_ram_read,
 -- Registers
 t8,
 n8,
 result,
 device_out_result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_return_output,
 device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_return_output,
 n8_MUX_uxn_opcodes_h_l502_c2_1228_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_return_output,
 result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_return_output,
 result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_return_output,
 t8_MUX_uxn_opcodes_h_l502_c2_1228_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_return_output,
 device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_return_output,
 n8_MUX_uxn_opcodes_h_l509_c7_95b1_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_return_output,
 result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_return_output,
 result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_return_output,
 t8_MUX_uxn_opcodes_h_l509_c7_95b1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_return_output,
 device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_return_output,
 n8_MUX_uxn_opcodes_h_l512_c7_21e6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_return_output,
 result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_return_output,
 result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_return_output,
 t8_MUX_uxn_opcodes_h_l512_c7_21e6_return_output,
 sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l519_c9_614a_return_output,
 MUX_uxn_opcodes_h_l519_c9_1c10_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l520_c42_ad6a_return_output,
 device_out_uxn_opcodes_h_l520_c23_fa5d_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : unsigned(0 downto 0);
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_iftrue : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_iffalse : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_return_output : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l502_c2_1228_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l502_c2_1228_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l502_c2_1228_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l502_c2_1228_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_cond : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_iftrue : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_iffalse : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_return_output : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_cond : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l506_c3_40e0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l502_c2_1228_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l502_c2_1228_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l509_c7_95b1_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l502_c2_1228_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l502_c2_1228_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse : unsigned(0 downto 0);
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_return_output : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l512_c7_21e6_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_return_output : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l510_c3_3d70 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l509_c7_95b1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l512_c7_21e6_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l509_c7_95b1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_iffalse : unsigned(0 downto 0);
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse : device_out_result_t;
 variable VAR_device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l512_c7_21e6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_cond : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse : unsigned(0 downto 0);
 variable VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_cond : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l518_c3_9718 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l512_c7_21e6_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l519_c9_1c10_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l519_c9_614a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l519_c9_614a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l519_c9_614a_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l519_c9_1c10_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l519_c9_1c10_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l519_c9_1c10_return_output : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_device_address : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_value : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_phase : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l520_c42_ad6a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l520_c42_ad6a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l520_c42_ad6a_return_output : unsigned(7 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_return_output : device_out_result_t;
 variable VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l521_c32_f6de_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_device_out_result_t_device_ram_address_d41d_uxn_opcodes_h_l522_c31_dd6f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_device_out_result_t_u8_value_d41d_uxn_opcodes_h_l523_c21_a6f4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_device_out_result_t_u16_addr_d41d_uxn_opcodes_h_l524_c22_cedd_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_vram_write_d41d_uxn_opcodes_h_l525_c26_b98f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_device_out_result_t_vram_write_layer_d41d_uxn_opcodes_h_l526_c29_5bd1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d_uxn_opcodes_h_l527_c24_e032_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_4aae_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_b1c2_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_2b1d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_1ed3_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_ec2b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_e09d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l509_l502_DUPLICATE_e449_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l509_l512_DUPLICATE_f706_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_23b1_uxn_opcodes_h_l530_l497_DUPLICATE_80c6_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
variable REG_VAR_device_out_result : device_out_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
  REG_VAR_device_out_result := device_out_result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l506_c3_40e0 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l506_c3_40e0;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l520_c42_ad6a_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_iftrue := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_y := resize(to_signed(-2, 3), 4);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l510_c3_3d70 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l510_c3_3d70;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l519_c9_614a_right := to_unsigned(3, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l518_c3_9718 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse := VAR_result_sp_relative_shift_uxn_opcodes_h_l518_c3_9718;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_device_ram_read := previous_device_ram_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse := VAR_CLOCK_ENABLE;
     VAR_device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_iftrue := device_out_result;
     VAR_device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue := device_out_result;
     VAR_device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue := device_out_result;
     VAR_sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_ins := VAR_ins;
     VAR_MUX_uxn_opcodes_h_l519_c9_1c10_iffalse := n8;
     VAR_n8_MUX_uxn_opcodes_h_l502_c2_1228_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l519_c9_614a_left := VAR_phase;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l520_c42_ad6a_left := VAR_phase;
     VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_previous_device_ram_read := VAR_previous_device_ram_read;
     VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_previous_ram_read := VAR_previous_ram_read;
     VAR_MUX_uxn_opcodes_h_l519_c9_1c10_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue := VAR_previous_stack_read;
     VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_device_address := t8;
     VAR_t8_MUX_uxn_opcodes_h_l502_c2_1228_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse := t8;
     -- sp_relative_shift[uxn_opcodes_h_l515_c30_e5ba] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_ins;
     sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_x <= VAR_sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_x;
     sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_y <= VAR_sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_return_output := sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l509_c7_95b1] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l509_c7_95b1_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_b1c2 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_b1c2_return_output := result.vram_write_layer;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_1ed3 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_1ed3_return_output := result.u16_value;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_4aae LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_4aae_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_e09d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_e09d_return_output := result.is_device_ram_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l509_l502_DUPLICATE_e449 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l509_l502_DUPLICATE_e449_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_2b1d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_2b1d_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l502_c6_d85c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_left;
     BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_return_output := BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_ec2b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_ec2b_return_output := result.device_ram_address;

     -- BIN_OP_EQ[uxn_opcodes_h_l512_c11_3193] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_left;
     BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_return_output := BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l509_l512_DUPLICATE_f706 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l509_l512_DUPLICATE_f706_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l519_c9_614a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l519_c9_614a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l519_c9_614a_left;
     BIN_OP_EQ_uxn_opcodes_h_l519_c9_614a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l519_c9_614a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l519_c9_614a_return_output := BIN_OP_EQ_uxn_opcodes_h_l519_c9_614a_return_output;

     -- BIN_OP_MINUS[uxn_opcodes_h_l520_c42_ad6a] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l520_c42_ad6a_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l520_c42_ad6a_left;
     BIN_OP_MINUS_uxn_opcodes_h_l520_c42_ad6a_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l520_c42_ad6a_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l520_c42_ad6a_return_output := BIN_OP_MINUS_uxn_opcodes_h_l520_c42_ad6a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l509_c11_500d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_left;
     BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_return_output := BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_return_output;

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l502_c2_1228_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l502_c2_1228_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l502_c6_d85c_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l509_c7_95b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l509_c7_95b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l509_c11_500d_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l512_c7_21e6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l512_c7_21e6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l512_c11_3193_return_output;
     VAR_MUX_uxn_opcodes_h_l519_c9_1c10_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l519_c9_614a_return_output;
     VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_phase := VAR_BIN_OP_MINUS_uxn_opcodes_h_l520_c42_ad6a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l509_l502_DUPLICATE_e449_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l509_l502_DUPLICATE_e449_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_1ed3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_1ed3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_1ed3_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_e09d_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_e09d_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_e09d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l509_l512_DUPLICATE_f706_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l509_l512_DUPLICATE_f706_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_2b1d_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_2b1d_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_2b1d_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_b1c2_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_b1c2_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_vram_write_layer_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_b1c2_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_ec2b_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_ec2b_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_ec2b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_4aae_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_4aae_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l509_l512_l502_DUPLICATE_4aae_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l509_c7_95b1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l515_c30_e5ba_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l509_c7_95b1] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l509_c7_95b1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l512_c7_21e6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_return_output;

     -- MUX[uxn_opcodes_h_l519_c9_1c10] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l519_c9_1c10_cond <= VAR_MUX_uxn_opcodes_h_l519_c9_1c10_cond;
     MUX_uxn_opcodes_h_l519_c9_1c10_iftrue <= VAR_MUX_uxn_opcodes_h_l519_c9_1c10_iftrue;
     MUX_uxn_opcodes_h_l519_c9_1c10_iffalse <= VAR_MUX_uxn_opcodes_h_l519_c9_1c10_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l519_c9_1c10_return_output := MUX_uxn_opcodes_h_l519_c9_1c10_return_output;

     -- t8_MUX[uxn_opcodes_h_l512_c7_21e6] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l512_c7_21e6_cond <= VAR_t8_MUX_uxn_opcodes_h_l512_c7_21e6_cond;
     t8_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue;
     t8_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l512_c7_21e6_return_output := t8_MUX_uxn_opcodes_h_l512_c7_21e6_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;
     VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_value := VAR_MUX_uxn_opcodes_h_l519_c9_1c10_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse := VAR_MUX_uxn_opcodes_h_l519_c9_1c10_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l512_c7_21e6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse := VAR_t8_MUX_uxn_opcodes_h_l512_c7_21e6_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l512_c7_21e6] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_return_output;

     -- t8_MUX[uxn_opcodes_h_l509_c7_95b1] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l509_c7_95b1_cond <= VAR_t8_MUX_uxn_opcodes_h_l509_c7_95b1_cond;
     t8_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue;
     t8_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l509_c7_95b1_return_output := t8_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;

     -- n8_MUX[uxn_opcodes_h_l512_c7_21e6] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l512_c7_21e6_cond <= VAR_n8_MUX_uxn_opcodes_h_l512_c7_21e6_cond;
     n8_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue;
     n8_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l512_c7_21e6_return_output := n8_MUX_uxn_opcodes_h_l512_c7_21e6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l509_c7_95b1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l502_c2_1228] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_return_output;

     -- Submodule level 3
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l512_c7_21e6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse := VAR_n8_MUX_uxn_opcodes_h_l512_c7_21e6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l502_c2_1228_iffalse := VAR_t8_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l517_c1_4eeb] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_return_output;

     -- t8_MUX[uxn_opcodes_h_l502_c2_1228] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l502_c2_1228_cond <= VAR_t8_MUX_uxn_opcodes_h_l502_c2_1228_cond;
     t8_MUX_uxn_opcodes_h_l502_c2_1228_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l502_c2_1228_iftrue;
     t8_MUX_uxn_opcodes_h_l502_c2_1228_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l502_c2_1228_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l502_c2_1228_return_output := t8_MUX_uxn_opcodes_h_l502_c2_1228_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l502_c2_1228] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_return_output;

     -- n8_MUX[uxn_opcodes_h_l509_c7_95b1] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l509_c7_95b1_cond <= VAR_n8_MUX_uxn_opcodes_h_l509_c7_95b1_cond;
     n8_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue;
     n8_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l509_c7_95b1_return_output := n8_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;

     -- Submodule level 4
     VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_CLOCK_ENABLE := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l517_c1_4eeb_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l502_c2_1228_iffalse := VAR_n8_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l502_c2_1228_return_output;
     -- device_out[uxn_opcodes_h_l520_c23_fa5d] LATENCY=0
     -- Clock enable
     device_out_uxn_opcodes_h_l520_c23_fa5d_CLOCK_ENABLE <= VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_CLOCK_ENABLE;
     -- Inputs
     device_out_uxn_opcodes_h_l520_c23_fa5d_device_address <= VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_device_address;
     device_out_uxn_opcodes_h_l520_c23_fa5d_value <= VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_value;
     device_out_uxn_opcodes_h_l520_c23_fa5d_phase <= VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_phase;
     device_out_uxn_opcodes_h_l520_c23_fa5d_previous_device_ram_read <= VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_previous_device_ram_read;
     device_out_uxn_opcodes_h_l520_c23_fa5d_previous_ram_read <= VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_previous_ram_read;
     -- Outputs
     VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_return_output := device_out_uxn_opcodes_h_l520_c23_fa5d_return_output;

     -- n8_MUX[uxn_opcodes_h_l502_c2_1228] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l502_c2_1228_cond <= VAR_n8_MUX_uxn_opcodes_h_l502_c2_1228_cond;
     n8_MUX_uxn_opcodes_h_l502_c2_1228_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l502_c2_1228_iftrue;
     n8_MUX_uxn_opcodes_h_l502_c2_1228_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l502_c2_1228_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l502_c2_1228_return_output := n8_MUX_uxn_opcodes_h_l502_c2_1228_return_output;

     -- Submodule level 5
     VAR_device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse := VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_return_output;
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l502_c2_1228_return_output;
     -- CONST_REF_RD_uint16_t_device_out_result_t_u16_addr_d41d[uxn_opcodes_h_l524_c22_cedd] LATENCY=0
     VAR_CONST_REF_RD_uint16_t_device_out_result_t_u16_addr_d41d_uxn_opcodes_h_l524_c22_cedd_return_output := VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_return_output.u16_addr;

     -- device_out_result_MUX[uxn_opcodes_h_l512_c7_21e6] LATENCY=0
     -- Inputs
     device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_cond <= VAR_device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_cond;
     device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue <= VAR_device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue;
     device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse <= VAR_device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse;
     -- Outputs
     VAR_device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_return_output := device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_return_output;

     -- CONST_REF_RD_uint1_t_device_out_result_t_vram_write_layer_d41d[uxn_opcodes_h_l526_c29_5bd1] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_out_result_t_vram_write_layer_d41d_uxn_opcodes_h_l526_c29_5bd1_return_output := VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_return_output.vram_write_layer;

     -- CONST_REF_RD_uint1_t_device_out_result_t_is_device_ram_write_d41d[uxn_opcodes_h_l521_c32_f6de] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l521_c32_f6de_return_output := VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_return_output.is_device_ram_write;

     -- CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d[uxn_opcodes_h_l527_c24_e032] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d_uxn_opcodes_h_l527_c24_e032_return_output := VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_return_output.is_deo_done;

     -- CONST_REF_RD_uint8_t_device_out_result_t_u8_value_d41d[uxn_opcodes_h_l523_c21_a6f4] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_out_result_t_u8_value_d41d_uxn_opcodes_h_l523_c21_a6f4_return_output := VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_return_output.u8_value;

     -- CONST_REF_RD_uint8_t_device_out_result_t_device_ram_address_d41d[uxn_opcodes_h_l522_c31_dd6f] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_out_result_t_device_ram_address_d41d_uxn_opcodes_h_l522_c31_dd6f_return_output := VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_return_output.device_ram_address;

     -- CONST_REF_RD_uint1_t_device_out_result_t_is_vram_write_d41d[uxn_opcodes_h_l525_c26_b98f] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_vram_write_d41d_uxn_opcodes_h_l525_c26_b98f_return_output := VAR_device_out_uxn_opcodes_h_l520_c23_fa5d_return_output.is_vram_write;

     -- Submodule level 6
     VAR_result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse := VAR_CONST_REF_RD_uint16_t_device_out_result_t_u16_addr_d41d_uxn_opcodes_h_l524_c22_cedd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse := VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_deo_done_d41d_uxn_opcodes_h_l527_c24_e032_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse := VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l521_c32_f6de_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse := VAR_CONST_REF_RD_uint1_t_device_out_result_t_is_vram_write_d41d_uxn_opcodes_h_l525_c26_b98f_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse := VAR_CONST_REF_RD_uint1_t_device_out_result_t_vram_write_layer_d41d_uxn_opcodes_h_l526_c29_5bd1_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse := VAR_CONST_REF_RD_uint8_t_device_out_result_t_device_ram_address_d41d_uxn_opcodes_h_l522_c31_dd6f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse := VAR_CONST_REF_RD_uint8_t_device_out_result_t_u8_value_d41d_uxn_opcodes_h_l523_c21_a6f4_return_output;
     VAR_device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse := VAR_device_out_result_MUX_uxn_opcodes_h_l512_c7_21e6_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l512_c7_21e6] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_cond;
     result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_return_output := result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l512_c7_21e6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_return_output := result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_return_output;

     -- result_is_device_ram_write_MUX[uxn_opcodes_h_l512_c7_21e6] LATENCY=0
     -- Inputs
     result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_cond <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_cond;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse;
     -- Outputs
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_return_output := result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l512_c7_21e6] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l512_c7_21e6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_return_output;

     -- result_device_ram_address_MUX[uxn_opcodes_h_l512_c7_21e6] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_return_output;

     -- device_out_result_MUX[uxn_opcodes_h_l509_c7_95b1] LATENCY=0
     -- Inputs
     device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_cond <= VAR_device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_cond;
     device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue <= VAR_device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue;
     device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse <= VAR_device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse;
     -- Outputs
     VAR_device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_return_output := device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;

     -- result_vram_write_layer_MUX[uxn_opcodes_h_l512_c7_21e6] LATENCY=0
     -- Inputs
     result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_cond <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_cond;
     result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_iftrue;
     result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_iffalse;
     -- Outputs
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_return_output := result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_return_output;

     -- Submodule level 7
     VAR_device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_iffalse := VAR_device_out_result_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l512_c7_21e6_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse := VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l512_c7_21e6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l512_c7_21e6_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse := VAR_result_is_vram_write_MUX_uxn_opcodes_h_l512_c7_21e6_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l512_c7_21e6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l512_c7_21e6_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse := VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l512_c7_21e6_return_output;
     -- result_is_device_ram_write_MUX[uxn_opcodes_h_l509_c7_95b1] LATENCY=0
     -- Inputs
     result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_cond <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_cond;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse;
     -- Outputs
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_return_output := result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;

     -- result_vram_write_layer_MUX[uxn_opcodes_h_l509_c7_95b1] LATENCY=0
     -- Inputs
     result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_cond <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_cond;
     result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue;
     result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse;
     -- Outputs
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_return_output := result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l509_c7_95b1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;

     -- device_out_result_MUX[uxn_opcodes_h_l502_c2_1228] LATENCY=0
     -- Inputs
     device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_cond <= VAR_device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_cond;
     device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_iftrue <= VAR_device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_iftrue;
     device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_iffalse <= VAR_device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_iffalse;
     -- Outputs
     VAR_device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_return_output := device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l509_c7_95b1] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;

     -- result_device_ram_address_MUX[uxn_opcodes_h_l509_c7_95b1] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l509_c7_95b1] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_cond;
     result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_return_output := result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l509_c7_95b1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_return_output := result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;

     -- Submodule level 8
     REG_VAR_device_out_result := VAR_device_out_result_MUX_uxn_opcodes_h_l502_c2_1228_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_iffalse := VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_iffalse := VAR_result_is_vram_write_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_iffalse := VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l509_c7_95b1_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l502_c2_1228] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_cond;
     result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_return_output := result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l502_c2_1228] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_return_output;

     -- result_is_device_ram_write_MUX[uxn_opcodes_h_l502_c2_1228] LATENCY=0
     -- Inputs
     result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_cond <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_cond;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_iftrue <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_iftrue;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_iffalse <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_iffalse;
     -- Outputs
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_return_output := result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_return_output;

     -- result_vram_write_layer_MUX[uxn_opcodes_h_l502_c2_1228] LATENCY=0
     -- Inputs
     result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_cond <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_cond;
     result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_iftrue <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_iftrue;
     result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_iffalse <= VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_iffalse;
     -- Outputs
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_return_output := result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l502_c2_1228] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_cond;
     result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_return_output := result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l502_c2_1228] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_return_output;

     -- result_device_ram_address_MUX[uxn_opcodes_h_l502_c2_1228] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_return_output;

     -- Submodule level 9
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_23b1_uxn_opcodes_h_l530_l497_DUPLICATE_80c6 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_23b1_uxn_opcodes_h_l530_l497_DUPLICATE_80c6_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_23b1(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l502_c2_1228_return_output,
     VAR_result_vram_write_layer_MUX_uxn_opcodes_h_l502_c2_1228_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l502_c2_1228_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l502_c2_1228_return_output,
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l502_c2_1228_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l502_c2_1228_return_output,
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l502_c2_1228_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l502_c2_1228_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l502_c2_1228_return_output);

     -- Submodule level 10
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_23b1_uxn_opcodes_h_l530_l497_DUPLICATE_80c6_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_23b1_uxn_opcodes_h_l530_l497_DUPLICATE_80c6_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
REG_COMB_device_out_result <= REG_VAR_device_out_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
     device_out_result <= REG_COMB_device_out_result;
 end if;
 end if;
end process;

end arch;
