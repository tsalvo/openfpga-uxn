-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity rot_0CLK_b288bfb7 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end rot_0CLK_b288bfb7;
architecture arch of rot_0CLK_b288bfb7 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal l8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_l8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2639_c6_04e9]
signal BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2639_c2_5a5d]
signal n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l2639_c2_5a5d]
signal l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2639_c2_5a5d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2639_c2_5a5d]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2639_c2_5a5d]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2639_c2_5a5d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2639_c2_5a5d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2639_c2_5a5d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2639_c2_5a5d]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2639_c2_5a5d]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2639_c2_5a5d]
signal result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2639_c2_5a5d]
signal t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2652_c11_a088]
signal BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2652_c7_c17b]
signal n8_MUX_uxn_opcodes_h_l2652_c7_c17b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l2652_c7_c17b]
signal l8_MUX_uxn_opcodes_h_l2652_c7_c17b_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2652_c7_c17b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2652_c7_c17b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2652_c7_c17b]
signal result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2652_c7_c17b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2652_c7_c17b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2652_c7_c17b]
signal t8_MUX_uxn_opcodes_h_l2652_c7_c17b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2655_c11_1f30]
signal BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2655_c7_e9c6]
signal n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l2655_c7_e9c6]
signal l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2655_c7_e9c6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2655_c7_e9c6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2655_c7_e9c6]
signal result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2655_c7_e9c6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2655_c7_e9c6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2655_c7_e9c6]
signal t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2659_c11_0ead]
signal BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2659_c7_4fb6]
signal n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l2659_c7_4fb6]
signal l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2659_c7_4fb6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2659_c7_4fb6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2659_c7_4fb6]
signal result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2659_c7_4fb6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2659_c7_4fb6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2661_c30_09b5]
signal sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2666_c11_10c1]
signal BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2666_c7_4215]
signal l8_MUX_uxn_opcodes_h_l2666_c7_4215_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2666_c7_4215_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2666_c7_4215]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2666_c7_4215]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2666_c7_4215]
signal result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2666_c7_4215]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2672_c11_a760]
signal BIN_OP_EQ_uxn_opcodes_h_l2672_c11_a760_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2672_c11_a760_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2672_c11_a760_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2672_c7_4edc]
signal result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2672_c7_4edc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2672_c7_4edc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8b52( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_opc_done := ref_toks_6;
      base.is_ram_write := ref_toks_7;
      base.is_vram_write := ref_toks_8;
      base.u8_value := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9
BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_left,
BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_right,
BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_return_output);

-- n8_MUX_uxn_opcodes_h_l2639_c2_5a5d
n8_MUX_uxn_opcodes_h_l2639_c2_5a5d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond,
n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue,
n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse,
n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output);

-- l8_MUX_uxn_opcodes_h_l2639_c2_5a5d
l8_MUX_uxn_opcodes_h_l2639_c2_5a5d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond,
l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue,
l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse,
l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond,
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output);

-- t8_MUX_uxn_opcodes_h_l2639_c2_5a5d
t8_MUX_uxn_opcodes_h_l2639_c2_5a5d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond,
t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue,
t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse,
t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088
BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_left,
BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_right,
BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_return_output);

-- n8_MUX_uxn_opcodes_h_l2652_c7_c17b
n8_MUX_uxn_opcodes_h_l2652_c7_c17b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2652_c7_c17b_cond,
n8_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue,
n8_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse,
n8_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output);

-- l8_MUX_uxn_opcodes_h_l2652_c7_c17b
l8_MUX_uxn_opcodes_h_l2652_c7_c17b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2652_c7_c17b_cond,
l8_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue,
l8_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse,
l8_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_cond,
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output);

-- t8_MUX_uxn_opcodes_h_l2652_c7_c17b
t8_MUX_uxn_opcodes_h_l2652_c7_c17b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2652_c7_c17b_cond,
t8_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue,
t8_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse,
t8_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30
BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_left,
BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_right,
BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_return_output);

-- n8_MUX_uxn_opcodes_h_l2655_c7_e9c6
n8_MUX_uxn_opcodes_h_l2655_c7_e9c6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond,
n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue,
n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse,
n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output);

-- l8_MUX_uxn_opcodes_h_l2655_c7_e9c6
l8_MUX_uxn_opcodes_h_l2655_c7_e9c6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond,
l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue,
l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse,
l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond,
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output);

-- t8_MUX_uxn_opcodes_h_l2655_c7_e9c6
t8_MUX_uxn_opcodes_h_l2655_c7_e9c6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond,
t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue,
t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse,
t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead
BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_left,
BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_right,
BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_return_output);

-- n8_MUX_uxn_opcodes_h_l2659_c7_4fb6
n8_MUX_uxn_opcodes_h_l2659_c7_4fb6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond,
n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue,
n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse,
n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output);

-- l8_MUX_uxn_opcodes_h_l2659_c7_4fb6
l8_MUX_uxn_opcodes_h_l2659_c7_4fb6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond,
l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue,
l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse,
l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond,
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5
sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_ins,
sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_x,
sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_y,
sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1
BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1_left,
BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1_right,
BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1_return_output);

-- l8_MUX_uxn_opcodes_h_l2666_c7_4215
l8_MUX_uxn_opcodes_h_l2666_c7_4215 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2666_c7_4215_cond,
l8_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue,
l8_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse,
l8_MUX_uxn_opcodes_h_l2666_c7_4215_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_cond,
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2672_c11_a760
BIN_OP_EQ_uxn_opcodes_h_l2672_c11_a760 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2672_c11_a760_left,
BIN_OP_EQ_uxn_opcodes_h_l2672_c11_a760_right,
BIN_OP_EQ_uxn_opcodes_h_l2672_c11_a760_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_cond,
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 l8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_return_output,
 n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output,
 l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output,
 t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_return_output,
 n8_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output,
 l8_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output,
 t8_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_return_output,
 n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output,
 l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output,
 t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_return_output,
 n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output,
 l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output,
 sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1_return_output,
 l8_MUX_uxn_opcodes_h_l2666_c7_4215_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2672_c11_a760_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2644_c3_2c9d : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2649_c3_d859 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2652_c7_c17b_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2652_c7_c17b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2653_c3_413a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2652_c7_c17b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2656_c3_8f11 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2666_c7_4215_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2663_c3_e8ca : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2666_c7_4215_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2669_c3_7cd4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2668_c3_cfc6 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_a760_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_a760_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_a760_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2673_c3_5931 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2672_c7_4edc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2652_l2655_l2672_l2639_DUPLICATE_4b94_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2652_l2666_l2655_DUPLICATE_c32c_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2659_l2652_l2655_DUPLICATE_7bb3_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2652_l2672_l2666_l2659_l2655_DUPLICATE_7553_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2678_l2635_DUPLICATE_2317_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_l8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_l8 := l8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2673_c3_5931 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2673_c3_5931;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2663_c3_e8ca := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2663_c3_e8ca;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2644_c3_2c9d := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2644_c3_2c9d;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_a760_right := to_unsigned(5, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2649_c3_d859 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2649_c3_d859;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2668_c3_cfc6 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2668_c3_cfc6;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_iftrue := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2656_c3_8f11 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2656_c3_8f11;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2669_c3_7cd4 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2669_c3_7cd4;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2653_c3_413a := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2653_c3_413a;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_ins := VAR_ins;
     VAR_l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse := l8;
     VAR_n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_a760_left := VAR_phase;
     VAR_l8_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse := t8;
     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2672_c7_4edc] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2672_c7_4edc_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2655_c11_1f30] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_left;
     BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_return_output := BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2639_c6_04e9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_left;
     BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_return_output := BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2659_l2652_l2655_DUPLICATE_7bb3 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2659_l2652_l2655_DUPLICATE_7bb3_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2666_c11_10c1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1_left;
     BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1_return_output := BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2661_c30_09b5] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_ins;
     sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_x;
     sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_return_output := sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2652_l2655_l2672_l2639_DUPLICATE_4b94 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2652_l2655_l2672_l2639_DUPLICATE_4b94_return_output := result.u8_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2652_l2666_l2655_DUPLICATE_c32c LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2652_l2666_l2655_DUPLICATE_c32c_return_output := result.sp_relative_shift;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2639_c2_5a5d] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2639_c2_5a5d_return_output := result.is_stack_index_flipped;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2639_c2_5a5d] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2639_c2_5a5d_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l2659_c11_0ead] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_left;
     BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_return_output := BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2652_l2672_l2666_l2659_l2655_DUPLICATE_7553 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2652_l2672_l2666_l2659_l2655_DUPLICATE_7553_return_output := result.is_opc_done;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2639_c2_5a5d] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2639_c2_5a5d_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2652_c11_a088] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_left;
     BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_return_output := BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2639_c2_5a5d] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2639_c2_5a5d_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2672_c11_a760] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2672_c11_a760_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_a760_left;
     BIN_OP_EQ_uxn_opcodes_h_l2672_c11_a760_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_a760_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_a760_return_output := BIN_OP_EQ_uxn_opcodes_h_l2672_c11_a760_return_output;

     -- Submodule level 1
     VAR_l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_04e9_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2652_c7_c17b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2652_c7_c17b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2652_c7_c17b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a088_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_1f30_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_0ead_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2666_c7_4215_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_10c1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_a760_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_a760_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_a760_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2652_l2666_l2655_DUPLICATE_c32c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2652_l2666_l2655_DUPLICATE_c32c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2652_l2666_l2655_DUPLICATE_c32c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2652_l2672_l2666_l2659_l2655_DUPLICATE_7553_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2652_l2672_l2666_l2659_l2655_DUPLICATE_7553_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2652_l2672_l2666_l2659_l2655_DUPLICATE_7553_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2652_l2672_l2666_l2659_l2655_DUPLICATE_7553_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2652_l2672_l2666_l2659_l2655_DUPLICATE_7553_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2659_l2652_l2655_DUPLICATE_7bb3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2659_l2652_l2655_DUPLICATE_7bb3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2659_l2652_l2655_DUPLICATE_7bb3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2652_l2655_l2672_l2639_DUPLICATE_4b94_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2652_l2655_l2672_l2639_DUPLICATE_4b94_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2652_l2655_l2672_l2639_DUPLICATE_4b94_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2652_l2655_l2672_l2639_DUPLICATE_4b94_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2639_c2_5a5d_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2639_c2_5a5d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2639_c2_5a5d_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2639_c2_5a5d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2672_c7_4edc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_09b5_return_output;
     -- n8_MUX[uxn_opcodes_h_l2659_c7_4fb6] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond <= VAR_n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond;
     n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue;
     n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output := n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2639_c2_5a5d] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2639_c2_5a5d] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2639_c2_5a5d] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2672_c7_4edc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_return_output;

     -- t8_MUX[uxn_opcodes_h_l2655_c7_e9c6] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond <= VAR_t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond;
     t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue;
     t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output := t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output;

     -- l8_MUX[uxn_opcodes_h_l2666_c7_4215] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2666_c7_4215_cond <= VAR_l8_MUX_uxn_opcodes_h_l2666_c7_4215_cond;
     l8_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue;
     l8_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2666_c7_4215_return_output := l8_MUX_uxn_opcodes_h_l2666_c7_4215_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2672_c7_4edc] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_return_output := result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2666_c7_4215] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2659_c7_4fb6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2639_c2_5a5d] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2672_c7_4edc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_return_output;

     -- Submodule level 2
     VAR_l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2666_c7_4215_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_4edc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_4215_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_4edc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_4edc_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output;
     -- l8_MUX[uxn_opcodes_h_l2659_c7_4fb6] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond <= VAR_l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond;
     l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue;
     l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output := l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2659_c7_4fb6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2655_c7_e9c6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2666_c7_4215] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_return_output := result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_return_output;

     -- n8_MUX[uxn_opcodes_h_l2655_c7_e9c6] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond <= VAR_n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond;
     n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue;
     n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output := n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2666_c7_4215] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_return_output;

     -- t8_MUX[uxn_opcodes_h_l2652_c7_c17b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2652_c7_c17b_cond <= VAR_t8_MUX_uxn_opcodes_h_l2652_c7_c17b_cond;
     t8_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue;
     t8_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output := t8_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2666_c7_4215] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_return_output;

     -- Submodule level 3
     VAR_l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_4215_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_4215_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_4215_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2652_c7_c17b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2659_c7_4fb6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output;

     -- l8_MUX[uxn_opcodes_h_l2655_c7_e9c6] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond <= VAR_l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond;
     l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue;
     l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output := l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output;

     -- t8_MUX[uxn_opcodes_h_l2639_c2_5a5d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond <= VAR_t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond;
     t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue;
     t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output := t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output;

     -- n8_MUX[uxn_opcodes_h_l2652_c7_c17b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2652_c7_c17b_cond <= VAR_n8_MUX_uxn_opcodes_h_l2652_c7_c17b_cond;
     n8_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue;
     n8_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output := n8_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2659_c7_4fb6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output := result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2655_c7_e9c6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2659_c7_4fb6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output;

     -- Submodule level 4
     VAR_l8_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_4fb6_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2655_c7_e9c6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2655_c7_e9c6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output;

     -- l8_MUX[uxn_opcodes_h_l2652_c7_c17b] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2652_c7_c17b_cond <= VAR_l8_MUX_uxn_opcodes_h_l2652_c7_c17b_cond;
     l8_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue;
     l8_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output := l8_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2639_c2_5a5d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2655_c7_e9c6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output := result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output;

     -- n8_MUX[uxn_opcodes_h_l2639_c2_5a5d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond <= VAR_n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond;
     n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue;
     n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output := n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2652_c7_c17b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output;

     -- Submodule level 5
     VAR_l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output;
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_e9c6_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2652_c7_c17b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2639_c2_5a5d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output;

     -- l8_MUX[uxn_opcodes_h_l2639_c2_5a5d] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond <= VAR_l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond;
     l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue;
     l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output := l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2652_c7_c17b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2652_c7_c17b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output := result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output;

     -- Submodule level 6
     REG_VAR_l8 := VAR_l8_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_c17b_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2639_c2_5a5d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2639_c2_5a5d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2639_c2_5a5d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output := result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2678_l2635_DUPLICATE_2317 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2678_l2635_DUPLICATE_2317_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8b52(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_5a5d_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2678_l2635_DUPLICATE_2317_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l2678_l2635_DUPLICATE_2317_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_l8 <= REG_VAR_l8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     l8 <= REG_COMB_l8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
