-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 52
entity jmp2_0CLK_9101a1df is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jmp2_0CLK_9101a1df;
architecture arch of jmp2_0CLK_9101a1df is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l656_c6_14dc]
signal BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l656_c1_b274]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l656_c2_83fe]
signal t16_MUX_uxn_opcodes_h_l656_c2_83fe_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l656_c2_83fe_return_output : unsigned(15 downto 0);

-- result_pc_MUX[uxn_opcodes_h_l656_c2_83fe]
signal result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_cond : unsigned(0 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_return_output : unsigned(15 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l656_c2_83fe]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l656_c2_83fe]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l656_c2_83fe]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_return_output : signed(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l656_c2_83fe]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l656_c2_83fe]
signal result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l657_c3_e6b0[uxn_opcodes_h_l657_c3_e6b0]
signal printf_uxn_opcodes_h_l657_c3_e6b0_uxn_opcodes_h_l657_c3_e6b0_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l661_c11_6031]
signal BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l661_c7_04db]
signal t16_MUX_uxn_opcodes_h_l661_c7_04db_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l661_c7_04db_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l661_c7_04db_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l661_c7_04db_return_output : unsigned(15 downto 0);

-- result_pc_MUX[uxn_opcodes_h_l661_c7_04db]
signal result_pc_MUX_uxn_opcodes_h_l661_c7_04db_cond : unsigned(0 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l661_c7_04db_iftrue : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l661_c7_04db_iffalse : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l661_c7_04db_return_output : unsigned(15 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l661_c7_04db]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l661_c7_04db]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l661_c7_04db]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_return_output : signed(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l661_c7_04db]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l661_c7_04db]
signal result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l664_c11_3a1a]
signal BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l664_c7_936f]
signal t16_MUX_uxn_opcodes_h_l664_c7_936f_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l664_c7_936f_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l664_c7_936f_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l664_c7_936f_return_output : unsigned(15 downto 0);

-- result_pc_MUX[uxn_opcodes_h_l664_c7_936f]
signal result_pc_MUX_uxn_opcodes_h_l664_c7_936f_cond : unsigned(0 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l664_c7_936f_iftrue : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l664_c7_936f_iffalse : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l664_c7_936f_return_output : unsigned(15 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l664_c7_936f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l664_c7_936f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l664_c7_936f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_return_output : signed(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l664_c7_936f]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l664_c7_936f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_return_output : unsigned(0 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l666_c3_d19d]
signal CONST_SL_8_uxn_opcodes_h_l666_c3_d19d_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l666_c3_d19d_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l669_c11_4f73]
signal BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l669_c7_bad3]
signal t16_MUX_uxn_opcodes_h_l669_c7_bad3_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l669_c7_bad3_return_output : unsigned(15 downto 0);

-- result_pc_MUX[uxn_opcodes_h_l669_c7_bad3]
signal result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_cond : unsigned(0 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_return_output : unsigned(15 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l669_c7_bad3]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l669_c7_bad3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l669_c7_bad3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_return_output : signed(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l669_c7_bad3]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l669_c7_bad3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l672_c11_4f91]
signal BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l672_c7_e3db]
signal t16_MUX_uxn_opcodes_h_l672_c7_e3db_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l672_c7_e3db_return_output : unsigned(15 downto 0);

-- result_pc_MUX[uxn_opcodes_h_l672_c7_e3db]
signal result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_cond : unsigned(0 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_return_output : unsigned(15 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l672_c7_e3db]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l672_c7_e3db]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_return_output : signed(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l672_c7_e3db]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l672_c7_e3db]
signal result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_return_output : unsigned(0 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l673_c3_dd6d]
signal BIN_OP_OR_uxn_opcodes_h_l673_c3_dd6d_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l673_c3_dd6d_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l673_c3_dd6d_return_output : unsigned(15 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l675_c32_4708]
signal BIN_OP_AND_uxn_opcodes_h_l675_c32_4708_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l675_c32_4708_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l675_c32_4708_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l675_c32_88cb]
signal BIN_OP_GT_uxn_opcodes_h_l675_c32_88cb_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l675_c32_88cb_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l675_c32_88cb_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l675_c32_9140]
signal MUX_uxn_opcodes_h_l675_c32_9140_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l675_c32_9140_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l675_c32_9140_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l675_c32_9140_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l679_c11_4206]
signal BIN_OP_EQ_uxn_opcodes_h_l679_c11_4206_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l679_c11_4206_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l679_c11_4206_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l679_c7_8cd4]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l679_c7_8cd4]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l679_c7_8cd4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_return_output : unsigned(0 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_f87d( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.pc := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.is_pc_updated := ref_toks_5;
      base.is_opc_done := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc
BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_left,
BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_right,
BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_return_output);

-- t16_MUX_uxn_opcodes_h_l656_c2_83fe
t16_MUX_uxn_opcodes_h_l656_c2_83fe : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l656_c2_83fe_cond,
t16_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue,
t16_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse,
t16_MUX_uxn_opcodes_h_l656_c2_83fe_return_output);

-- result_pc_MUX_uxn_opcodes_h_l656_c2_83fe
result_pc_MUX_uxn_opcodes_h_l656_c2_83fe : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_cond,
result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue,
result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse,
result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe
result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe
result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe
result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe
result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_return_output);

-- printf_uxn_opcodes_h_l657_c3_e6b0_uxn_opcodes_h_l657_c3_e6b0
printf_uxn_opcodes_h_l657_c3_e6b0_uxn_opcodes_h_l657_c3_e6b0 : entity work.printf_uxn_opcodes_h_l657_c3_e6b0_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l657_c3_e6b0_uxn_opcodes_h_l657_c3_e6b0_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031
BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_left,
BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_right,
BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_return_output);

-- t16_MUX_uxn_opcodes_h_l661_c7_04db
t16_MUX_uxn_opcodes_h_l661_c7_04db : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l661_c7_04db_cond,
t16_MUX_uxn_opcodes_h_l661_c7_04db_iftrue,
t16_MUX_uxn_opcodes_h_l661_c7_04db_iffalse,
t16_MUX_uxn_opcodes_h_l661_c7_04db_return_output);

-- result_pc_MUX_uxn_opcodes_h_l661_c7_04db
result_pc_MUX_uxn_opcodes_h_l661_c7_04db : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_pc_MUX_uxn_opcodes_h_l661_c7_04db_cond,
result_pc_MUX_uxn_opcodes_h_l661_c7_04db_iftrue,
result_pc_MUX_uxn_opcodes_h_l661_c7_04db_iffalse,
result_pc_MUX_uxn_opcodes_h_l661_c7_04db_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db
result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db
result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db
result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db
result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a
BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_left,
BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_right,
BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_return_output);

-- t16_MUX_uxn_opcodes_h_l664_c7_936f
t16_MUX_uxn_opcodes_h_l664_c7_936f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l664_c7_936f_cond,
t16_MUX_uxn_opcodes_h_l664_c7_936f_iftrue,
t16_MUX_uxn_opcodes_h_l664_c7_936f_iffalse,
t16_MUX_uxn_opcodes_h_l664_c7_936f_return_output);

-- result_pc_MUX_uxn_opcodes_h_l664_c7_936f
result_pc_MUX_uxn_opcodes_h_l664_c7_936f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_pc_MUX_uxn_opcodes_h_l664_c7_936f_cond,
result_pc_MUX_uxn_opcodes_h_l664_c7_936f_iftrue,
result_pc_MUX_uxn_opcodes_h_l664_c7_936f_iffalse,
result_pc_MUX_uxn_opcodes_h_l664_c7_936f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f
result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f
result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f
result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f
result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_return_output);

-- CONST_SL_8_uxn_opcodes_h_l666_c3_d19d
CONST_SL_8_uxn_opcodes_h_l666_c3_d19d : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l666_c3_d19d_x,
CONST_SL_8_uxn_opcodes_h_l666_c3_d19d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73
BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_left,
BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_right,
BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_return_output);

-- t16_MUX_uxn_opcodes_h_l669_c7_bad3
t16_MUX_uxn_opcodes_h_l669_c7_bad3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l669_c7_bad3_cond,
t16_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue,
t16_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse,
t16_MUX_uxn_opcodes_h_l669_c7_bad3_return_output);

-- result_pc_MUX_uxn_opcodes_h_l669_c7_bad3
result_pc_MUX_uxn_opcodes_h_l669_c7_bad3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_cond,
result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue,
result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse,
result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3
result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3
result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3
result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3
result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91
BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91_left,
BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91_right,
BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91_return_output);

-- t16_MUX_uxn_opcodes_h_l672_c7_e3db
t16_MUX_uxn_opcodes_h_l672_c7_e3db : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l672_c7_e3db_cond,
t16_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue,
t16_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse,
t16_MUX_uxn_opcodes_h_l672_c7_e3db_return_output);

-- result_pc_MUX_uxn_opcodes_h_l672_c7_e3db
result_pc_MUX_uxn_opcodes_h_l672_c7_e3db : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_cond,
result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue,
result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse,
result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db
result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db
result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db
result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db
result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l673_c3_dd6d
BIN_OP_OR_uxn_opcodes_h_l673_c3_dd6d : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l673_c3_dd6d_left,
BIN_OP_OR_uxn_opcodes_h_l673_c3_dd6d_right,
BIN_OP_OR_uxn_opcodes_h_l673_c3_dd6d_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l675_c32_4708
BIN_OP_AND_uxn_opcodes_h_l675_c32_4708 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l675_c32_4708_left,
BIN_OP_AND_uxn_opcodes_h_l675_c32_4708_right,
BIN_OP_AND_uxn_opcodes_h_l675_c32_4708_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l675_c32_88cb
BIN_OP_GT_uxn_opcodes_h_l675_c32_88cb : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l675_c32_88cb_left,
BIN_OP_GT_uxn_opcodes_h_l675_c32_88cb_right,
BIN_OP_GT_uxn_opcodes_h_l675_c32_88cb_return_output);

-- MUX_uxn_opcodes_h_l675_c32_9140
MUX_uxn_opcodes_h_l675_c32_9140 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l675_c32_9140_cond,
MUX_uxn_opcodes_h_l675_c32_9140_iftrue,
MUX_uxn_opcodes_h_l675_c32_9140_iffalse,
MUX_uxn_opcodes_h_l675_c32_9140_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l679_c11_4206
BIN_OP_EQ_uxn_opcodes_h_l679_c11_4206 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l679_c11_4206_left,
BIN_OP_EQ_uxn_opcodes_h_l679_c11_4206_right,
BIN_OP_EQ_uxn_opcodes_h_l679_c11_4206_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4
result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4
result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4
result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_return_output,
 t16_MUX_uxn_opcodes_h_l656_c2_83fe_return_output,
 result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_return_output,
 t16_MUX_uxn_opcodes_h_l661_c7_04db_return_output,
 result_pc_MUX_uxn_opcodes_h_l661_c7_04db_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_return_output,
 t16_MUX_uxn_opcodes_h_l664_c7_936f_return_output,
 result_pc_MUX_uxn_opcodes_h_l664_c7_936f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_return_output,
 CONST_SL_8_uxn_opcodes_h_l666_c3_d19d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_return_output,
 t16_MUX_uxn_opcodes_h_l669_c7_bad3_return_output,
 result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91_return_output,
 t16_MUX_uxn_opcodes_h_l672_c7_e3db_return_output,
 result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_return_output,
 BIN_OP_OR_uxn_opcodes_h_l673_c3_dd6d_return_output,
 BIN_OP_AND_uxn_opcodes_h_l675_c32_4708_return_output,
 BIN_OP_GT_uxn_opcodes_h_l675_c32_88cb_return_output,
 MUX_uxn_opcodes_h_l675_c32_9140_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l679_c11_4206_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_iffalse : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l661_c7_04db_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l656_c2_83fe_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l656_c2_83fe_cond : unsigned(0 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l661_c7_04db_return_output : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_return_output : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l658_c3_75b5 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l657_c3_e6b0_uxn_opcodes_h_l657_c3_e6b0_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l661_c7_04db_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l661_c7_04db_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l664_c7_936f_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l661_c7_04db_cond : unsigned(0 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l661_c7_04db_iftrue : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l661_c7_04db_iffalse : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l664_c7_936f_return_output : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l661_c7_04db_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l662_c3_d129 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l664_c7_936f_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l664_c7_936f_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l669_c7_bad3_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l664_c7_936f_cond : unsigned(0 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l664_c7_936f_iftrue : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l664_c7_936f_iffalse : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_return_output : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l664_c7_936f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l667_c3_99d4 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l666_c3_d19d_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l666_c3_d19d_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l672_c7_e3db_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l669_c7_bad3_cond : unsigned(0 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_return_output : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l670_c3_d731 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l669_c7_bad3_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l672_c7_e3db_cond : unsigned(0 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l673_c3_dd6d_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l673_c3_dd6d_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l673_c3_dd6d_return_output : unsigned(15 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l675_c32_9140_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l675_c32_9140_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l675_c32_9140_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l675_c32_4708_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l675_c32_4708_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l675_c32_4708_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l675_c32_88cb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l675_c32_88cb_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l675_c32_88cb_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l675_c32_9140_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l679_c11_4206_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l679_c11_4206_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l679_c11_4206_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l669_l656_l672_l661_l664_DUPLICATE_3833_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l669_l656_l661_l679_l664_DUPLICATE_c5f3_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l669_l656_l672_l661_l664_DUPLICATE_d54a_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l669_l656_l661_l679_l664_DUPLICATE_2d2e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l669_l672_l661_l679_l664_DUPLICATE_0bf5_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l665_l673_DUPLICATE_3562_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_f87d_uxn_opcodes_h_l685_l652_DUPLICATE_3638_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l658_c3_75b5 := resize(to_unsigned(2, 2), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l658_c3_75b5;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91_right := to_unsigned(4, 3);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l667_c3_99d4 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l667_c3_99d4;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l662_c3_d129 := resize(to_unsigned(2, 2), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l662_c3_d129;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l670_c3_d731 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l670_c3_d731;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_right := to_unsigned(3, 2);
     VAR_BIN_OP_AND_uxn_opcodes_h_l675_c32_4708_right := to_unsigned(128, 8);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_right := to_unsigned(2, 2);
     VAR_MUX_uxn_opcodes_h_l675_c32_9140_iftrue := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_MUX_uxn_opcodes_h_l675_c32_9140_iffalse := resize(to_signed(-2, 3), 8);
     VAR_BIN_OP_GT_uxn_opcodes_h_l675_c32_88cb_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l679_c11_4206_right := to_unsigned(5, 3);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_AND_uxn_opcodes_h_l675_c32_4708_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l679_c11_4206_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l673_c3_dd6d_left := t16;
     VAR_t16_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l661_c7_04db_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse := t16;
     -- CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l669_l656_l672_l661_l664_DUPLICATE_3833 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l669_l656_l672_l661_l664_DUPLICATE_3833_return_output := result.pc;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l669_l656_l672_l661_l664_DUPLICATE_d54a LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l669_l656_l672_l661_l664_DUPLICATE_d54a_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l661_c11_6031] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_left;
     BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_return_output := BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l669_l656_l661_l679_l664_DUPLICATE_2d2e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l669_l656_l661_l679_l664_DUPLICATE_2d2e_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l664_c11_3a1a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_left;
     BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_return_output := BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l672_c11_4f91] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91_left;
     BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91_return_output := BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l679_c11_4206] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l679_c11_4206_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l679_c11_4206_left;
     BIN_OP_EQ_uxn_opcodes_h_l679_c11_4206_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l679_c11_4206_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l679_c11_4206_return_output := BIN_OP_EQ_uxn_opcodes_h_l679_c11_4206_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l656_c6_14dc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_left;
     BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_return_output := BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l669_l656_l661_l679_l664_DUPLICATE_c5f3 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l669_l656_l661_l679_l664_DUPLICATE_c5f3_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l669_c11_4f73] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_left;
     BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_return_output := BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_return_output;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l665_l673_DUPLICATE_3562 LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l665_l673_DUPLICATE_3562_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l669_l672_l661_l679_l664_DUPLICATE_0bf5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l669_l672_l661_l679_l664_DUPLICATE_0bf5_return_output := result.is_opc_done;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l669_c7_bad3] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l669_c7_bad3_return_output := result.stack_address_sp_offset;

     -- BIN_OP_AND[uxn_opcodes_h_l675_c32_4708] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l675_c32_4708_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l675_c32_4708_left;
     BIN_OP_AND_uxn_opcodes_h_l675_c32_4708_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l675_c32_4708_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l675_c32_4708_return_output := BIN_OP_AND_uxn_opcodes_h_l675_c32_4708_return_output;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l675_c32_88cb_left := VAR_BIN_OP_AND_uxn_opcodes_h_l675_c32_4708_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l656_c2_83fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l656_c6_14dc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l661_c7_04db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l661_c7_04db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_6031_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l664_c7_936f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l664_c7_936f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l664_c11_3a1a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l669_c7_bad3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l669_c11_4f73_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l672_c7_e3db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l672_c11_4f91_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l679_c11_4206_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l679_c11_4206_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l679_c11_4206_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l673_c3_dd6d_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l665_l673_DUPLICATE_3562_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l666_c3_d19d_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l665_l673_DUPLICATE_3562_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l669_l656_l672_l661_l664_DUPLICATE_d54a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l669_l656_l672_l661_l664_DUPLICATE_d54a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l669_l656_l672_l661_l664_DUPLICATE_d54a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l669_l656_l672_l661_l664_DUPLICATE_d54a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l669_l656_l672_l661_l664_DUPLICATE_d54a_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l669_l656_l672_l661_l664_DUPLICATE_3833_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l661_c7_04db_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l669_l656_l672_l661_l664_DUPLICATE_3833_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l664_c7_936f_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l669_l656_l672_l661_l664_DUPLICATE_3833_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l669_l656_l672_l661_l664_DUPLICATE_3833_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l669_l656_l672_l661_l664_DUPLICATE_3833_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l669_l672_l661_l679_l664_DUPLICATE_0bf5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l669_l672_l661_l679_l664_DUPLICATE_0bf5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l669_l672_l661_l679_l664_DUPLICATE_0bf5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l669_l672_l661_l679_l664_DUPLICATE_0bf5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l669_l672_l661_l679_l664_DUPLICATE_0bf5_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l669_l656_l661_l679_l664_DUPLICATE_2d2e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l669_l656_l661_l679_l664_DUPLICATE_2d2e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l669_l656_l661_l679_l664_DUPLICATE_2d2e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l669_l656_l661_l679_l664_DUPLICATE_2d2e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l669_l656_l661_l679_l664_DUPLICATE_2d2e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l669_l656_l661_l679_l664_DUPLICATE_c5f3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l669_l656_l661_l679_l664_DUPLICATE_c5f3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l669_l656_l661_l679_l664_DUPLICATE_c5f3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l669_l656_l661_l679_l664_DUPLICATE_c5f3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l669_l656_l661_l679_l664_DUPLICATE_c5f3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l669_c7_bad3_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l669_c7_bad3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l679_c7_8cd4] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l679_c7_8cd4] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l673_c3_dd6d] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l673_c3_dd6d_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l673_c3_dd6d_left;
     BIN_OP_OR_uxn_opcodes_h_l673_c3_dd6d_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l673_c3_dd6d_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l673_c3_dd6d_return_output := BIN_OP_OR_uxn_opcodes_h_l673_c3_dd6d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l679_c7_8cd4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l675_c32_88cb] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l675_c32_88cb_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l675_c32_88cb_left;
     BIN_OP_GT_uxn_opcodes_h_l675_c32_88cb_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l675_c32_88cb_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l675_c32_88cb_return_output := BIN_OP_GT_uxn_opcodes_h_l675_c32_88cb_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l666_c3_d19d] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l666_c3_d19d_x <= VAR_CONST_SL_8_uxn_opcodes_h_l666_c3_d19d_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l666_c3_d19d_return_output := CONST_SL_8_uxn_opcodes_h_l666_c3_d19d_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l656_c1_b274] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l675_c32_9140_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l675_c32_88cb_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l673_c3_dd6d_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l673_c3_dd6d_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l664_c7_936f_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l666_c3_d19d_return_output;
     VAR_printf_uxn_opcodes_h_l657_c3_e6b0_uxn_opcodes_h_l657_c3_e6b0_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l656_c1_b274_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l679_c7_8cd4_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l679_c7_8cd4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l679_c7_8cd4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l669_c7_bad3_return_output;
     -- printf_uxn_opcodes_h_l657_c3_e6b0[uxn_opcodes_h_l657_c3_e6b0] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l657_c3_e6b0_uxn_opcodes_h_l657_c3_e6b0_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l657_c3_e6b0_uxn_opcodes_h_l657_c3_e6b0_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- t16_MUX[uxn_opcodes_h_l672_c7_e3db] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l672_c7_e3db_cond <= VAR_t16_MUX_uxn_opcodes_h_l672_c7_e3db_cond;
     t16_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue;
     t16_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l672_c7_e3db_return_output := t16_MUX_uxn_opcodes_h_l672_c7_e3db_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l672_c7_e3db] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l672_c7_e3db] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_return_output;

     -- MUX[uxn_opcodes_h_l675_c32_9140] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l675_c32_9140_cond <= VAR_MUX_uxn_opcodes_h_l675_c32_9140_cond;
     MUX_uxn_opcodes_h_l675_c32_9140_iftrue <= VAR_MUX_uxn_opcodes_h_l675_c32_9140_iftrue;
     MUX_uxn_opcodes_h_l675_c32_9140_iffalse <= VAR_MUX_uxn_opcodes_h_l675_c32_9140_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l675_c32_9140_return_output := MUX_uxn_opcodes_h_l675_c32_9140_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l664_c7_936f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l672_c7_e3db] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_return_output;

     -- result_pc_MUX[uxn_opcodes_h_l672_c7_e3db] LATENCY=0
     -- Inputs
     result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_cond <= VAR_result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_cond;
     result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue <= VAR_result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue;
     result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse <= VAR_result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse;
     -- Outputs
     VAR_result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_return_output := result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue := VAR_MUX_uxn_opcodes_h_l675_c32_9140_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l672_c7_e3db_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l672_c7_e3db_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l672_c7_e3db_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse := VAR_result_pc_MUX_uxn_opcodes_h_l672_c7_e3db_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l664_c7_936f_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse := VAR_t16_MUX_uxn_opcodes_h_l672_c7_e3db_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l672_c7_e3db] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l661_c7_04db] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l669_c7_bad3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l669_c7_bad3] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l669_c7_bad3] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_return_output;

     -- result_pc_MUX[uxn_opcodes_h_l669_c7_bad3] LATENCY=0
     -- Inputs
     result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_cond <= VAR_result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_cond;
     result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue <= VAR_result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue;
     result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse <= VAR_result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse;
     -- Outputs
     VAR_result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_return_output := result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_return_output;

     -- t16_MUX[uxn_opcodes_h_l669_c7_bad3] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l669_c7_bad3_cond <= VAR_t16_MUX_uxn_opcodes_h_l669_c7_bad3_cond;
     t16_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue;
     t16_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l669_c7_bad3_return_output := t16_MUX_uxn_opcodes_h_l669_c7_bad3_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l669_c7_bad3_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l669_c7_bad3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l669_c7_bad3_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l664_c7_936f_iffalse := VAR_result_pc_MUX_uxn_opcodes_h_l669_c7_bad3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l672_c7_e3db_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l661_c7_04db_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l664_c7_936f_iffalse := VAR_t16_MUX_uxn_opcodes_h_l669_c7_bad3_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l656_c2_83fe] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l664_c7_936f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_return_output;

     -- result_pc_MUX[uxn_opcodes_h_l664_c7_936f] LATENCY=0
     -- Inputs
     result_pc_MUX_uxn_opcodes_h_l664_c7_936f_cond <= VAR_result_pc_MUX_uxn_opcodes_h_l664_c7_936f_cond;
     result_pc_MUX_uxn_opcodes_h_l664_c7_936f_iftrue <= VAR_result_pc_MUX_uxn_opcodes_h_l664_c7_936f_iftrue;
     result_pc_MUX_uxn_opcodes_h_l664_c7_936f_iffalse <= VAR_result_pc_MUX_uxn_opcodes_h_l664_c7_936f_iffalse;
     -- Outputs
     VAR_result_pc_MUX_uxn_opcodes_h_l664_c7_936f_return_output := result_pc_MUX_uxn_opcodes_h_l664_c7_936f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l664_c7_936f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l669_c7_bad3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l664_c7_936f] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_return_output;

     -- t16_MUX[uxn_opcodes_h_l664_c7_936f] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l664_c7_936f_cond <= VAR_t16_MUX_uxn_opcodes_h_l664_c7_936f_cond;
     t16_MUX_uxn_opcodes_h_l664_c7_936f_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l664_c7_936f_iftrue;
     t16_MUX_uxn_opcodes_h_l664_c7_936f_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l664_c7_936f_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l664_c7_936f_return_output := t16_MUX_uxn_opcodes_h_l664_c7_936f_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l664_c7_936f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l664_c7_936f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l664_c7_936f_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l661_c7_04db_iffalse := VAR_result_pc_MUX_uxn_opcodes_h_l664_c7_936f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l669_c7_bad3_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l661_c7_04db_iffalse := VAR_t16_MUX_uxn_opcodes_h_l664_c7_936f_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l664_c7_936f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l661_c7_04db] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l661_c7_04db] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l661_c7_04db] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_return_output;

     -- t16_MUX[uxn_opcodes_h_l661_c7_04db] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l661_c7_04db_cond <= VAR_t16_MUX_uxn_opcodes_h_l661_c7_04db_cond;
     t16_MUX_uxn_opcodes_h_l661_c7_04db_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l661_c7_04db_iftrue;
     t16_MUX_uxn_opcodes_h_l661_c7_04db_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l661_c7_04db_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l661_c7_04db_return_output := t16_MUX_uxn_opcodes_h_l661_c7_04db_return_output;

     -- result_pc_MUX[uxn_opcodes_h_l661_c7_04db] LATENCY=0
     -- Inputs
     result_pc_MUX_uxn_opcodes_h_l661_c7_04db_cond <= VAR_result_pc_MUX_uxn_opcodes_h_l661_c7_04db_cond;
     result_pc_MUX_uxn_opcodes_h_l661_c7_04db_iftrue <= VAR_result_pc_MUX_uxn_opcodes_h_l661_c7_04db_iftrue;
     result_pc_MUX_uxn_opcodes_h_l661_c7_04db_iffalse <= VAR_result_pc_MUX_uxn_opcodes_h_l661_c7_04db_iffalse;
     -- Outputs
     VAR_result_pc_MUX_uxn_opcodes_h_l661_c7_04db_return_output := result_pc_MUX_uxn_opcodes_h_l661_c7_04db_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_04db_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_04db_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l661_c7_04db_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse := VAR_result_pc_MUX_uxn_opcodes_h_l661_c7_04db_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l664_c7_936f_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse := VAR_t16_MUX_uxn_opcodes_h_l661_c7_04db_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l656_c2_83fe] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_return_output;

     -- t16_MUX[uxn_opcodes_h_l656_c2_83fe] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l656_c2_83fe_cond <= VAR_t16_MUX_uxn_opcodes_h_l656_c2_83fe_cond;
     t16_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue;
     t16_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l656_c2_83fe_return_output := t16_MUX_uxn_opcodes_h_l656_c2_83fe_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l661_c7_04db] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l656_c2_83fe] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l656_c2_83fe] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_return_output;

     -- result_pc_MUX[uxn_opcodes_h_l656_c2_83fe] LATENCY=0
     -- Inputs
     result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_cond <= VAR_result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_cond;
     result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue <= VAR_result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue;
     result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse <= VAR_result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse;
     -- Outputs
     VAR_result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_return_output := result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_return_output;

     -- Submodule level 7
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_04db_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l656_c2_83fe_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l656_c2_83fe] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_return_output;

     -- Submodule level 8
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_f87d_uxn_opcodes_h_l685_l652_DUPLICATE_3638 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_f87d_uxn_opcodes_h_l685_l652_DUPLICATE_3638_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_f87d(
     result,
     VAR_result_pc_MUX_uxn_opcodes_h_l656_c2_83fe_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l656_c2_83fe_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l656_c2_83fe_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l656_c2_83fe_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l656_c2_83fe_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l656_c2_83fe_return_output);

     -- Submodule level 9
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_f87d_uxn_opcodes_h_l685_l652_DUPLICATE_3638_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_f87d_uxn_opcodes_h_l685_l652_DUPLICATE_3638_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
