-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 54
entity div_0CLK_af9273cc is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end div_0CLK_af9273cc;
architecture arch of div_0CLK_af9273cc is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2185_c6_44cb]
signal BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2185_c1_2a50]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2185_c2_aa93]
signal n8_MUX_uxn_opcodes_h_l2185_c2_aa93_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2185_c2_aa93]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2185_c2_aa93]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2185_c2_aa93]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2185_c2_aa93]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2185_c2_aa93]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2185_c2_aa93]
signal result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2185_c2_aa93]
signal t8_MUX_uxn_opcodes_h_l2185_c2_aa93_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l2186_c3_e09e[uxn_opcodes_h_l2186_c3_e09e]
signal printf_uxn_opcodes_h_l2186_c3_e09e_uxn_opcodes_h_l2186_c3_e09e_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2190_c11_dd2d]
signal BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2190_c7_b4a9]
signal n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2190_c7_b4a9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2190_c7_b4a9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2190_c7_b4a9]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2190_c7_b4a9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2190_c7_b4a9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2190_c7_b4a9]
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2190_c7_b4a9]
signal t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2193_c11_7fd2]
signal BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2193_c7_4b62]
signal n8_MUX_uxn_opcodes_h_l2193_c7_4b62_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2193_c7_4b62]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2193_c7_4b62]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2193_c7_4b62]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2193_c7_4b62]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2193_c7_4b62]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2193_c7_4b62]
signal result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2193_c7_4b62]
signal t8_MUX_uxn_opcodes_h_l2193_c7_4b62_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2197_c11_36fa]
signal BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2197_c7_0d1f]
signal n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2197_c7_0d1f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2197_c7_0d1f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2197_c7_0d1f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2197_c7_0d1f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2197_c7_0d1f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2197_c7_0d1f]
signal result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2200_c11_d6ab]
signal BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2200_c7_54e8]
signal n8_MUX_uxn_opcodes_h_l2200_c7_54e8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2200_c7_54e8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2200_c7_54e8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2200_c7_54e8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2200_c7_54e8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2200_c7_54e8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2200_c7_54e8]
signal result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2203_c30_773f]
signal sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2206_c21_0844]
signal BIN_OP_EQ_uxn_opcodes_h_l2206_c21_0844_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2206_c21_0844_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2206_c21_0844_return_output : unsigned(0 downto 0);

-- BIN_OP_DIV[uxn_opcodes_h_l2206_c35_a6c6]
signal BIN_OP_DIV_uxn_opcodes_h_l2206_c35_a6c6_left : unsigned(7 downto 0);
signal BIN_OP_DIV_uxn_opcodes_h_l2206_c35_a6c6_right : unsigned(7 downto 0);
signal BIN_OP_DIV_uxn_opcodes_h_l2206_c35_a6c6_return_output : unsigned(7 downto 0);

-- MUX[uxn_opcodes_h_l2206_c21_b71b]
signal MUX_uxn_opcodes_h_l2206_c21_b71b_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l2206_c21_b71b_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l2206_c21_b71b_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l2206_c21_b71b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2208_c11_b45d]
signal BIN_OP_EQ_uxn_opcodes_h_l2208_c11_b45d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2208_c11_b45d_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2208_c11_b45d_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2208_c7_acdd]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2208_c7_acdd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2208_c7_acdd]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8cda( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb
BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_left,
BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_right,
BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_return_output);

-- n8_MUX_uxn_opcodes_h_l2185_c2_aa93
n8_MUX_uxn_opcodes_h_l2185_c2_aa93 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2185_c2_aa93_cond,
n8_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue,
n8_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse,
n8_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93
result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93
result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93
result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93
result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93
result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_cond,
result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output);

-- t8_MUX_uxn_opcodes_h_l2185_c2_aa93
t8_MUX_uxn_opcodes_h_l2185_c2_aa93 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2185_c2_aa93_cond,
t8_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue,
t8_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse,
t8_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output);

-- printf_uxn_opcodes_h_l2186_c3_e09e_uxn_opcodes_h_l2186_c3_e09e
printf_uxn_opcodes_h_l2186_c3_e09e_uxn_opcodes_h_l2186_c3_e09e : entity work.printf_uxn_opcodes_h_l2186_c3_e09e_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2186_c3_e09e_uxn_opcodes_h_l2186_c3_e09e_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d
BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_left,
BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_right,
BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_return_output);

-- n8_MUX_uxn_opcodes_h_l2190_c7_b4a9
n8_MUX_uxn_opcodes_h_l2190_c7_b4a9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond,
n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue,
n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse,
n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9
result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond,
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output);

-- t8_MUX_uxn_opcodes_h_l2190_c7_b4a9
t8_MUX_uxn_opcodes_h_l2190_c7_b4a9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond,
t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue,
t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse,
t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2
BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_left,
BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_right,
BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_return_output);

-- n8_MUX_uxn_opcodes_h_l2193_c7_4b62
n8_MUX_uxn_opcodes_h_l2193_c7_4b62 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2193_c7_4b62_cond,
n8_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue,
n8_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse,
n8_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62
result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62
result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62
result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62
result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62
result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_cond,
result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output);

-- t8_MUX_uxn_opcodes_h_l2193_c7_4b62
t8_MUX_uxn_opcodes_h_l2193_c7_4b62 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2193_c7_4b62_cond,
t8_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue,
t8_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse,
t8_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa
BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_left,
BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_right,
BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_return_output);

-- n8_MUX_uxn_opcodes_h_l2197_c7_0d1f
n8_MUX_uxn_opcodes_h_l2197_c7_0d1f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond,
n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue,
n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse,
n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f
result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f
result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab
BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_left,
BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_right,
BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_return_output);

-- n8_MUX_uxn_opcodes_h_l2200_c7_54e8
n8_MUX_uxn_opcodes_h_l2200_c7_54e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2200_c7_54e8_cond,
n8_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue,
n8_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse,
n8_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8
result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8
result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8
result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8
result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8
result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_cond,
result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2203_c30_773f
sp_relative_shift_uxn_opcodes_h_l2203_c30_773f : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_ins,
sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_x,
sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_y,
sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2206_c21_0844
BIN_OP_EQ_uxn_opcodes_h_l2206_c21_0844 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2206_c21_0844_left,
BIN_OP_EQ_uxn_opcodes_h_l2206_c21_0844_right,
BIN_OP_EQ_uxn_opcodes_h_l2206_c21_0844_return_output);

-- BIN_OP_DIV_uxn_opcodes_h_l2206_c35_a6c6
BIN_OP_DIV_uxn_opcodes_h_l2206_c35_a6c6 : entity work.BIN_OP_DIV_uint8_t_uint8_t_0CLK_a148083c port map (
BIN_OP_DIV_uxn_opcodes_h_l2206_c35_a6c6_left,
BIN_OP_DIV_uxn_opcodes_h_l2206_c35_a6c6_right,
BIN_OP_DIV_uxn_opcodes_h_l2206_c35_a6c6_return_output);

-- MUX_uxn_opcodes_h_l2206_c21_b71b
MUX_uxn_opcodes_h_l2206_c21_b71b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l2206_c21_b71b_cond,
MUX_uxn_opcodes_h_l2206_c21_b71b_iftrue,
MUX_uxn_opcodes_h_l2206_c21_b71b_iffalse,
MUX_uxn_opcodes_h_l2206_c21_b71b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2208_c11_b45d
BIN_OP_EQ_uxn_opcodes_h_l2208_c11_b45d : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2208_c11_b45d_left,
BIN_OP_EQ_uxn_opcodes_h_l2208_c11_b45d_right,
BIN_OP_EQ_uxn_opcodes_h_l2208_c11_b45d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd
result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd
result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd
result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_return_output,
 n8_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output,
 t8_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_return_output,
 n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output,
 t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_return_output,
 n8_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output,
 t8_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_return_output,
 n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_return_output,
 n8_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output,
 sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2206_c21_0844_return_output,
 BIN_OP_DIV_uxn_opcodes_h_l2206_c35_a6c6_return_output,
 MUX_uxn_opcodes_h_l2206_c21_b71b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2208_c11_b45d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2185_c2_aa93_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2187_c3_1492 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2185_c2_aa93_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2186_c3_e09e_uxn_opcodes_h_l2186_c3_e09e_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2191_c3_388a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2193_c7_4b62_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2195_c3_d1da : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2193_c7_4b62_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2198_c3_1823 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2200_c7_54e8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2205_c3_35ca : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2200_c7_54e8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2206_c21_b71b_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2206_c21_b71b_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2206_c21_b71b_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2206_c21_0844_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2206_c21_0844_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2206_c21_0844_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l2206_c35_a6c6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l2206_c35_a6c6_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l2206_c35_a6c6_return_output : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2206_c21_b71b_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2208_c11_b45d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2208_c11_b45d_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2208_c11_b45d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2200_l2197_l2193_l2190_l2185_DUPLICATE_1ce8_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2208_l2197_l2193_l2190_l2185_DUPLICATE_f645_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2208_l2197_l2193_l2190_l2185_DUPLICATE_2aa8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2200_l2197_l2193_l2190_l2185_DUPLICATE_4c7f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2208_l2200_l2197_l2193_l2190_DUPLICATE_7905_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l2214_l2181_DUPLICATE_d0db_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2198_c3_1823 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2198_c3_1823;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2205_c3_35ca := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2205_c3_35ca;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2191_c3_388a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2191_c3_388a;
     VAR_sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2206_c21_0844_right := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2208_c11_b45d_right := to_unsigned(5, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2195_c3_d1da := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2195_c3_d1da;
     VAR_MUX_uxn_opcodes_h_l2206_c21_b71b_iftrue := resize(to_unsigned(0, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2187_c3_1492 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2187_c3_1492;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2208_c11_b45d_left := VAR_phase;
     VAR_BIN_OP_DIV_uxn_opcodes_h_l2206_c35_a6c6_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_DIV_uxn_opcodes_h_l2206_c35_a6c6_right := t8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2206_c21_0844_left := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse := t8;
     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2200_c7_54e8] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2200_c7_54e8_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2200_l2197_l2193_l2190_l2185_DUPLICATE_1ce8 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2200_l2197_l2193_l2190_l2185_DUPLICATE_1ce8_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2200_c11_d6ab] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_left;
     BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_return_output := BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2197_c11_36fa] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_left;
     BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_return_output := BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2203_c30_773f] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_ins;
     sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_x;
     sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_return_output := sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2208_l2197_l2193_l2190_l2185_DUPLICATE_2aa8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2208_l2197_l2193_l2190_l2185_DUPLICATE_2aa8_return_output := result.is_stack_write;

     -- BIN_OP_DIV[uxn_opcodes_h_l2206_c35_a6c6] LATENCY=0
     -- Inputs
     BIN_OP_DIV_uxn_opcodes_h_l2206_c35_a6c6_left <= VAR_BIN_OP_DIV_uxn_opcodes_h_l2206_c35_a6c6_left;
     BIN_OP_DIV_uxn_opcodes_h_l2206_c35_a6c6_right <= VAR_BIN_OP_DIV_uxn_opcodes_h_l2206_c35_a6c6_right;
     -- Outputs
     VAR_BIN_OP_DIV_uxn_opcodes_h_l2206_c35_a6c6_return_output := BIN_OP_DIV_uxn_opcodes_h_l2206_c35_a6c6_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2190_c11_dd2d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_left;
     BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_return_output := BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2206_c21_0844] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2206_c21_0844_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2206_c21_0844_left;
     BIN_OP_EQ_uxn_opcodes_h_l2206_c21_0844_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2206_c21_0844_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2206_c21_0844_return_output := BIN_OP_EQ_uxn_opcodes_h_l2206_c21_0844_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2200_l2197_l2193_l2190_l2185_DUPLICATE_4c7f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2200_l2197_l2193_l2190_l2185_DUPLICATE_4c7f_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2208_l2200_l2197_l2193_l2190_DUPLICATE_7905 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2208_l2200_l2197_l2193_l2190_DUPLICATE_7905_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2185_c6_44cb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_left;
     BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_return_output := BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2208_l2197_l2193_l2190_l2185_DUPLICATE_f645 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2208_l2197_l2193_l2190_l2185_DUPLICATE_f645_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2208_c11_b45d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2208_c11_b45d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2208_c11_b45d_left;
     BIN_OP_EQ_uxn_opcodes_h_l2208_c11_b45d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2208_c11_b45d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2208_c11_b45d_return_output := BIN_OP_EQ_uxn_opcodes_h_l2208_c11_b45d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2193_c11_7fd2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_left;
     BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_return_output := BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_return_output;

     -- Submodule level 1
     VAR_MUX_uxn_opcodes_h_l2206_c21_b71b_iffalse := VAR_BIN_OP_DIV_uxn_opcodes_h_l2206_c35_a6c6_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2185_c2_aa93_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2185_c2_aa93_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2185_c6_44cb_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_dd2d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2193_c7_4b62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2193_c7_4b62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2193_c11_7fd2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_36fa_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2200_c7_54e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_d6ab_return_output;
     VAR_MUX_uxn_opcodes_h_l2206_c21_b71b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2206_c21_0844_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2208_c11_b45d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2208_c11_b45d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2208_c11_b45d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2200_l2197_l2193_l2190_l2185_DUPLICATE_1ce8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2200_l2197_l2193_l2190_l2185_DUPLICATE_1ce8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2200_l2197_l2193_l2190_l2185_DUPLICATE_1ce8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2200_l2197_l2193_l2190_l2185_DUPLICATE_1ce8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2200_l2197_l2193_l2190_l2185_DUPLICATE_1ce8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2208_l2200_l2197_l2193_l2190_DUPLICATE_7905_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2208_l2200_l2197_l2193_l2190_DUPLICATE_7905_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2208_l2200_l2197_l2193_l2190_DUPLICATE_7905_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2208_l2200_l2197_l2193_l2190_DUPLICATE_7905_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2208_l2200_l2197_l2193_l2190_DUPLICATE_7905_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2208_l2197_l2193_l2190_l2185_DUPLICATE_f645_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2208_l2197_l2193_l2190_l2185_DUPLICATE_f645_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2208_l2197_l2193_l2190_l2185_DUPLICATE_f645_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2208_l2197_l2193_l2190_l2185_DUPLICATE_f645_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2208_l2197_l2193_l2190_l2185_DUPLICATE_f645_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2208_l2197_l2193_l2190_l2185_DUPLICATE_2aa8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2208_l2197_l2193_l2190_l2185_DUPLICATE_2aa8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2208_l2197_l2193_l2190_l2185_DUPLICATE_2aa8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2208_l2197_l2193_l2190_l2185_DUPLICATE_2aa8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2208_l2197_l2193_l2190_l2185_DUPLICATE_2aa8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2200_l2197_l2193_l2190_l2185_DUPLICATE_4c7f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2200_l2197_l2193_l2190_l2185_DUPLICATE_4c7f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2200_l2197_l2193_l2190_l2185_DUPLICATE_4c7f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2200_l2197_l2193_l2190_l2185_DUPLICATE_4c7f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2200_l2197_l2193_l2190_l2185_DUPLICATE_4c7f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2200_c7_54e8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2203_c30_773f_return_output;
     -- n8_MUX[uxn_opcodes_h_l2200_c7_54e8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2200_c7_54e8_cond <= VAR_n8_MUX_uxn_opcodes_h_l2200_c7_54e8_cond;
     n8_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue;
     n8_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output := n8_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2208_c7_acdd] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_return_output;

     -- t8_MUX[uxn_opcodes_h_l2193_c7_4b62] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2193_c7_4b62_cond <= VAR_t8_MUX_uxn_opcodes_h_l2193_c7_4b62_cond;
     t8_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue;
     t8_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output := t8_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2200_c7_54e8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2185_c1_2a50] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_return_output;

     -- MUX[uxn_opcodes_h_l2206_c21_b71b] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l2206_c21_b71b_cond <= VAR_MUX_uxn_opcodes_h_l2206_c21_b71b_cond;
     MUX_uxn_opcodes_h_l2206_c21_b71b_iftrue <= VAR_MUX_uxn_opcodes_h_l2206_c21_b71b_iftrue;
     MUX_uxn_opcodes_h_l2206_c21_b71b_iffalse <= VAR_MUX_uxn_opcodes_h_l2206_c21_b71b_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l2206_c21_b71b_return_output := MUX_uxn_opcodes_h_l2206_c21_b71b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2208_c7_acdd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2200_c7_54e8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2208_c7_acdd] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue := VAR_MUX_uxn_opcodes_h_l2206_c21_b71b_return_output;
     VAR_printf_uxn_opcodes_h_l2186_c3_e09e_uxn_opcodes_h_l2186_c3_e09e_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2185_c1_2a50_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2208_c7_acdd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2208_c7_acdd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2208_c7_acdd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2200_c7_54e8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2197_c7_0d1f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output;

     -- printf_uxn_opcodes_h_l2186_c3_e09e[uxn_opcodes_h_l2186_c3_e09e] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2186_c3_e09e_uxn_opcodes_h_l2186_c3_e09e_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2186_c3_e09e_uxn_opcodes_h_l2186_c3_e09e_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2197_c7_0d1f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output;

     -- t8_MUX[uxn_opcodes_h_l2190_c7_b4a9] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond <= VAR_t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond;
     t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue;
     t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output := t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2200_c7_54e8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output;

     -- n8_MUX[uxn_opcodes_h_l2197_c7_0d1f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond <= VAR_n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond;
     n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue;
     n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output := n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2200_c7_54e8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2200_c7_54e8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output := result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2200_c7_54e8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2197_c7_0d1f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output;

     -- t8_MUX[uxn_opcodes_h_l2185_c2_aa93] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2185_c2_aa93_cond <= VAR_t8_MUX_uxn_opcodes_h_l2185_c2_aa93_cond;
     t8_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue;
     t8_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output := t8_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output;

     -- n8_MUX[uxn_opcodes_h_l2193_c7_4b62] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2193_c7_4b62_cond <= VAR_n8_MUX_uxn_opcodes_h_l2193_c7_4b62_cond;
     n8_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue;
     n8_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output := n8_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2197_c7_0d1f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2197_c7_0d1f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2193_c7_4b62] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2197_c7_0d1f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2193_c7_4b62] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0d1f_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2193_c7_4b62] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output;

     -- n8_MUX[uxn_opcodes_h_l2190_c7_b4a9] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond <= VAR_n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond;
     n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue;
     n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output := n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2193_c7_4b62] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2193_c7_4b62] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output := result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2190_c7_b4a9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2190_c7_b4a9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2193_c7_4b62] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2193_c7_4b62_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2185_c2_aa93] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2190_c7_b4a9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output := result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output;

     -- n8_MUX[uxn_opcodes_h_l2185_c2_aa93] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2185_c2_aa93_cond <= VAR_n8_MUX_uxn_opcodes_h_l2185_c2_aa93_cond;
     n8_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue;
     n8_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output := n8_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2190_c7_b4a9] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2190_c7_b4a9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2190_c7_b4a9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2185_c2_aa93] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_b4a9_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2185_c2_aa93] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output := result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2185_c2_aa93] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2185_c2_aa93] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2185_c2_aa93] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l2214_l2181_DUPLICATE_d0db LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l2214_l2181_DUPLICATE_d0db_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8cda(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2185_c2_aa93_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l2214_l2181_DUPLICATE_d0db_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l2214_l2181_DUPLICATE_d0db_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
