-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity sta_0CLK_bce25fe8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sta_0CLK_bce25fe8;
architecture arch of sta_0CLK_bce25fe8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2298_c6_2afb]
signal BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2298_c2_0b27]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2298_c2_0b27]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2298_c2_0b27]
signal result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2298_c2_0b27]
signal result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2298_c2_0b27]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2298_c2_0b27]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2298_c2_0b27]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2298_c2_0b27]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2298_c2_0b27]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2298_c2_0b27]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2298_c2_0b27]
signal t16_MUX_uxn_opcodes_h_l2298_c2_0b27_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(15 downto 0);

-- n8_MUX[uxn_opcodes_h_l2298_c2_0b27]
signal n8_MUX_uxn_opcodes_h_l2298_c2_0b27_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2311_c11_35e4]
signal BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2311_c7_c001]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2311_c7_c001]
signal result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2311_c7_c001]
signal result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2311_c7_c001]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2311_c7_c001]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2311_c7_c001]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2311_c7_c001]
signal t16_MUX_uxn_opcodes_h_l2311_c7_c001_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2311_c7_c001_return_output : unsigned(15 downto 0);

-- n8_MUX[uxn_opcodes_h_l2311_c7_c001]
signal n8_MUX_uxn_opcodes_h_l2311_c7_c001_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2311_c7_c001_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2314_c11_3b19]
signal BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2314_c7_e15b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2314_c7_e15b]
signal result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2314_c7_e15b]
signal result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2314_c7_e15b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2314_c7_e15b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2314_c7_e15b]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2314_c7_e15b]
signal t16_MUX_uxn_opcodes_h_l2314_c7_e15b_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output : unsigned(15 downto 0);

-- n8_MUX[uxn_opcodes_h_l2314_c7_e15b]
signal n8_MUX_uxn_opcodes_h_l2314_c7_e15b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output : unsigned(7 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l2316_c3_a632]
signal CONST_SL_8_uxn_opcodes_h_l2316_c3_a632_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l2316_c3_a632_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2319_c11_1c0b]
signal BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2319_c7_c757]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2319_c7_c757]
signal result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2319_c7_c757]
signal result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2319_c7_c757]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2319_c7_c757]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2319_c7_c757]
signal t16_MUX_uxn_opcodes_h_l2319_c7_c757_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2319_c7_c757_return_output : unsigned(15 downto 0);

-- n8_MUX[uxn_opcodes_h_l2319_c7_c757]
signal n8_MUX_uxn_opcodes_h_l2319_c7_c757_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2319_c7_c757_return_output : unsigned(7 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l2320_c3_8dac]
signal BIN_OP_OR_uxn_opcodes_h_l2320_c3_8dac_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2320_c3_8dac_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2320_c3_8dac_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2322_c11_48e7]
signal BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2322_c7_aed6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2322_c7_aed6]
signal result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2322_c7_aed6]
signal result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2322_c7_aed6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2322_c7_aed6]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2322_c7_aed6]
signal n8_MUX_uxn_opcodes_h_l2322_c7_aed6_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2324_c30_04f9]
signal sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_return_output : signed(3 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_500b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_pc_updated := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.u16_value := ref_toks_4;
      base.is_ram_write := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_stack_write := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_stack_index_flipped := ref_toks_9;
      base.is_opc_done := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb
BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_left,
BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_right,
BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27
result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27
result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27
result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_cond,
result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27
result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_cond,
result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27
result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27
result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27
result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27
result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output);

-- t16_MUX_uxn_opcodes_h_l2298_c2_0b27
t16_MUX_uxn_opcodes_h_l2298_c2_0b27 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2298_c2_0b27_cond,
t16_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue,
t16_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse,
t16_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output);

-- n8_MUX_uxn_opcodes_h_l2298_c2_0b27
n8_MUX_uxn_opcodes_h_l2298_c2_0b27 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2298_c2_0b27_cond,
n8_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue,
n8_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse,
n8_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4
BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_left,
BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_right,
BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001
result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001
result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_cond,
result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001
result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_cond,
result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001
result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001
result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_return_output);

-- t16_MUX_uxn_opcodes_h_l2311_c7_c001
t16_MUX_uxn_opcodes_h_l2311_c7_c001 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2311_c7_c001_cond,
t16_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue,
t16_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse,
t16_MUX_uxn_opcodes_h_l2311_c7_c001_return_output);

-- n8_MUX_uxn_opcodes_h_l2311_c7_c001
n8_MUX_uxn_opcodes_h_l2311_c7_c001 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2311_c7_c001_cond,
n8_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue,
n8_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse,
n8_MUX_uxn_opcodes_h_l2311_c7_c001_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19
BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_left,
BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_right,
BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b
result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b
result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_cond,
result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b
result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_cond,
result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b
result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b
result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output);

-- t16_MUX_uxn_opcodes_h_l2314_c7_e15b
t16_MUX_uxn_opcodes_h_l2314_c7_e15b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2314_c7_e15b_cond,
t16_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue,
t16_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse,
t16_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output);

-- n8_MUX_uxn_opcodes_h_l2314_c7_e15b
n8_MUX_uxn_opcodes_h_l2314_c7_e15b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2314_c7_e15b_cond,
n8_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue,
n8_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse,
n8_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output);

-- CONST_SL_8_uxn_opcodes_h_l2316_c3_a632
CONST_SL_8_uxn_opcodes_h_l2316_c3_a632 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l2316_c3_a632_x,
CONST_SL_8_uxn_opcodes_h_l2316_c3_a632_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b
BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_left,
BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_right,
BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757
result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757
result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_cond,
result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757
result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_cond,
result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757
result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757
result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_return_output);

-- t16_MUX_uxn_opcodes_h_l2319_c7_c757
t16_MUX_uxn_opcodes_h_l2319_c7_c757 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2319_c7_c757_cond,
t16_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue,
t16_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse,
t16_MUX_uxn_opcodes_h_l2319_c7_c757_return_output);

-- n8_MUX_uxn_opcodes_h_l2319_c7_c757
n8_MUX_uxn_opcodes_h_l2319_c7_c757 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2319_c7_c757_cond,
n8_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue,
n8_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse,
n8_MUX_uxn_opcodes_h_l2319_c7_c757_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l2320_c3_8dac
BIN_OP_OR_uxn_opcodes_h_l2320_c3_8dac : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l2320_c3_8dac_left,
BIN_OP_OR_uxn_opcodes_h_l2320_c3_8dac_right,
BIN_OP_OR_uxn_opcodes_h_l2320_c3_8dac_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7
BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7_left,
BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7_right,
BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6
result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6
result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_cond,
result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6
result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_cond,
result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6
result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6
result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output);

-- n8_MUX_uxn_opcodes_h_l2322_c7_aed6
n8_MUX_uxn_opcodes_h_l2322_c7_aed6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2322_c7_aed6_cond,
n8_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue,
n8_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse,
n8_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9
sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_ins,
sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_x,
sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_y,
sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output,
 t16_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output,
 n8_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_return_output,
 t16_MUX_uxn_opcodes_h_l2311_c7_c001_return_output,
 n8_MUX_uxn_opcodes_h_l2311_c7_c001_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output,
 t16_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output,
 n8_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output,
 CONST_SL_8_uxn_opcodes_h_l2316_c3_a632_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_return_output,
 t16_MUX_uxn_opcodes_h_l2319_c7_c757_return_output,
 n8_MUX_uxn_opcodes_h_l2319_c7_c757_return_output,
 BIN_OP_OR_uxn_opcodes_h_l2320_c3_8dac_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output,
 n8_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output,
 sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2303_c3_63f6 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2308_c3_d686 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2311_c7_c001_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2298_c2_0b27_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2311_c7_c001_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2298_c2_0b27_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2312_c3_edcd : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2311_c7_c001_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2311_c7_c001_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2317_c3_c5a3 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2314_c7_e15b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2319_c7_c757_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2314_c7_e15b_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2319_c7_c757_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2314_c7_e15b_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2316_c3_a632_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2316_c3_a632_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2319_c7_c757_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2319_c7_c757_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2320_c3_8dac_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2320_c3_8dac_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2320_c3_8dac_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2322_c7_aed6_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2314_l2311_l2298_l2322_l2319_DUPLICATE_e800_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2314_l2311_l2298_l2322_l2319_DUPLICATE_1ce9_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2311_l2322_l2314_l2319_DUPLICATE_f77f_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2311_l2322_l2314_l2319_DUPLICATE_6706_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2311_l2322_l2314_l2319_DUPLICATE_663b_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2315_l2320_DUPLICATE_bf86_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_500b_uxn_opcodes_h_l2293_l2331_DUPLICATE_50a1_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2317_c3_c5a3 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2317_c3_c5a3;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_y := resize(to_signed(-3, 3), 4);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2303_c3_63f6 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2303_c3_63f6;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7_right := to_unsigned(4, 3);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2312_c3_edcd := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2312_c3_edcd;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2308_c3_d686 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2308_c3_d686;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2320_c3_8dac_left := t16;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse := t16;
     -- BIN_OP_EQ[uxn_opcodes_h_l2311_c11_35e4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_left;
     BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_return_output := BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_return_output;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2315_l2320_DUPLICATE_bf86 LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2315_l2320_DUPLICATE_bf86_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2311_l2322_l2314_l2319_DUPLICATE_663b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2311_l2322_l2314_l2319_DUPLICATE_663b_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2298_c6_2afb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_left;
     BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_return_output := BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2314_c7_e15b] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2314_c7_e15b_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2314_c11_3b19] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_left;
     BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_return_output := BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2319_c11_1c0b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_left;
     BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_return_output := BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2322_c11_48e7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7_left;
     BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7_return_output := BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2298_c2_0b27] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2298_c2_0b27_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2314_l2311_l2298_l2322_l2319_DUPLICATE_e800 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2314_l2311_l2298_l2322_l2319_DUPLICATE_e800_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2311_l2322_l2314_l2319_DUPLICATE_6706 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2311_l2322_l2314_l2319_DUPLICATE_6706_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2314_l2311_l2298_l2322_l2319_DUPLICATE_1ce9 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2314_l2311_l2298_l2322_l2319_DUPLICATE_1ce9_return_output := result.u16_value;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2298_c2_0b27] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2298_c2_0b27_return_output := result.is_vram_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2311_l2322_l2314_l2319_DUPLICATE_f77f LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2311_l2322_l2314_l2319_DUPLICATE_f77f_return_output := result.sp_relative_shift;

     -- result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d[uxn_opcodes_h_l2298_c2_0b27] LATENCY=0
     VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2298_c2_0b27_return_output := result.is_stack_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2298_c2_0b27] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2298_c2_0b27_return_output := result.is_pc_updated;

     -- sp_relative_shift[uxn_opcodes_h_l2324_c30_04f9] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_ins;
     sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_x;
     sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_return_output := sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l2298_c2_0b27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2298_c2_0b27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2298_c6_2afb_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2311_c7_c001_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2311_c7_c001_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2311_c11_35e4_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2314_c7_e15b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2314_c7_e15b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2314_c11_3b19_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2319_c7_c757_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2319_c7_c757_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2319_c11_1c0b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2322_c7_aed6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2322_c11_48e7_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2320_c3_8dac_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2315_l2320_DUPLICATE_bf86_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l2316_c3_a632_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2315_l2320_DUPLICATE_bf86_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2311_l2322_l2314_l2319_DUPLICATE_f77f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2311_l2322_l2314_l2319_DUPLICATE_f77f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2311_l2322_l2314_l2319_DUPLICATE_f77f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2311_l2322_l2314_l2319_DUPLICATE_f77f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2314_l2311_l2298_l2322_l2319_DUPLICATE_1ce9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2314_l2311_l2298_l2322_l2319_DUPLICATE_1ce9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2314_l2311_l2298_l2322_l2319_DUPLICATE_1ce9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2314_l2311_l2298_l2322_l2319_DUPLICATE_1ce9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2314_l2311_l2298_l2322_l2319_DUPLICATE_1ce9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2311_l2322_l2314_l2319_DUPLICATE_6706_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2311_l2322_l2314_l2319_DUPLICATE_6706_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2311_l2322_l2314_l2319_DUPLICATE_6706_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2311_l2322_l2314_l2319_DUPLICATE_6706_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2311_l2322_l2314_l2319_DUPLICATE_663b_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2311_l2322_l2314_l2319_DUPLICATE_663b_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2311_l2322_l2314_l2319_DUPLICATE_663b_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2311_l2322_l2314_l2319_DUPLICATE_663b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2314_l2311_l2298_l2322_l2319_DUPLICATE_e800_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2314_l2311_l2298_l2322_l2319_DUPLICATE_e800_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2314_l2311_l2298_l2322_l2319_DUPLICATE_e800_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2314_l2311_l2298_l2322_l2319_DUPLICATE_e800_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2314_l2311_l2298_l2322_l2319_DUPLICATE_e800_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2298_c2_0b27_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2298_c2_0b27_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse := VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2298_c2_0b27_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2298_c2_0b27_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2314_c7_e15b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2324_c30_04f9_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2314_c7_e15b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2322_c7_aed6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2322_c7_aed6] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output := result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l2316_c3_a632] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l2316_c3_a632_x <= VAR_CONST_SL_8_uxn_opcodes_h_l2316_c3_a632_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l2316_c3_a632_return_output := CONST_SL_8_uxn_opcodes_h_l2316_c3_a632_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2298_c2_0b27] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2298_c2_0b27] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2298_c2_0b27] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output;

     -- n8_MUX[uxn_opcodes_h_l2322_c7_aed6] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2322_c7_aed6_cond <= VAR_n8_MUX_uxn_opcodes_h_l2322_c7_aed6_cond;
     n8_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue;
     n8_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output := n8_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l2320_c3_8dac] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l2320_c3_8dac_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l2320_c3_8dac_left;
     BIN_OP_OR_uxn_opcodes_h_l2320_c3_8dac_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l2320_c3_8dac_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l2320_c3_8dac_return_output := BIN_OP_OR_uxn_opcodes_h_l2320_c3_8dac_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2322_c7_aed6] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2322_c7_aed6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2322_c7_aed6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output := result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2298_c2_0b27] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output;

     -- Submodule level 2
     VAR_t16_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l2320_c3_8dac_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l2316_c3_a632_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2322_c7_aed6_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2319_c7_c757] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_return_output;

     -- t16_MUX[uxn_opcodes_h_l2319_c7_c757] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2319_c7_c757_cond <= VAR_t16_MUX_uxn_opcodes_h_l2319_c7_c757_cond;
     t16_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue;
     t16_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2319_c7_c757_return_output := t16_MUX_uxn_opcodes_h_l2319_c7_c757_return_output;

     -- n8_MUX[uxn_opcodes_h_l2319_c7_c757] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2319_c7_c757_cond <= VAR_n8_MUX_uxn_opcodes_h_l2319_c7_c757_cond;
     n8_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue;
     n8_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2319_c7_c757_return_output := n8_MUX_uxn_opcodes_h_l2319_c7_c757_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2319_c7_c757] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2319_c7_c757] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2319_c7_c757] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_return_output := result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2311_c7_c001] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2319_c7_c757] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_return_output := result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2319_c7_c757_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2319_c7_c757_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2319_c7_c757_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2319_c7_c757_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2311_c7_c001_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2319_c7_c757_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2319_c7_c757_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2319_c7_c757_return_output;
     -- n8_MUX[uxn_opcodes_h_l2314_c7_e15b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2314_c7_e15b_cond <= VAR_n8_MUX_uxn_opcodes_h_l2314_c7_e15b_cond;
     n8_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue;
     n8_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output := n8_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2314_c7_e15b] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output;

     -- t16_MUX[uxn_opcodes_h_l2314_c7_e15b] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2314_c7_e15b_cond <= VAR_t16_MUX_uxn_opcodes_h_l2314_c7_e15b_cond;
     t16_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue;
     t16_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output := t16_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2314_c7_e15b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2314_c7_e15b] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output := result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2298_c2_0b27] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2314_c7_e15b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output := result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2314_c7_e15b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2314_c7_e15b_return_output;
     -- n8_MUX[uxn_opcodes_h_l2311_c7_c001] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2311_c7_c001_cond <= VAR_n8_MUX_uxn_opcodes_h_l2311_c7_c001_cond;
     n8_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue;
     n8_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2311_c7_c001_return_output := n8_MUX_uxn_opcodes_h_l2311_c7_c001_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2311_c7_c001] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_return_output := result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2311_c7_c001] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_return_output;

     -- t16_MUX[uxn_opcodes_h_l2311_c7_c001] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2311_c7_c001_cond <= VAR_t16_MUX_uxn_opcodes_h_l2311_c7_c001_cond;
     t16_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue;
     t16_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2311_c7_c001_return_output := t16_MUX_uxn_opcodes_h_l2311_c7_c001_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2311_c7_c001] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2311_c7_c001] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_return_output := result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2311_c7_c001] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2311_c7_c001_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2311_c7_c001_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2311_c7_c001_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2311_c7_c001_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2311_c7_c001_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2311_c7_c001_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2311_c7_c001_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2298_c2_0b27] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2298_c2_0b27] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output := result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output;

     -- n8_MUX[uxn_opcodes_h_l2298_c2_0b27] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2298_c2_0b27_cond <= VAR_n8_MUX_uxn_opcodes_h_l2298_c2_0b27_cond;
     n8_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue;
     n8_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output := n8_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2298_c2_0b27] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2298_c2_0b27] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output := result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output;

     -- t16_MUX[uxn_opcodes_h_l2298_c2_0b27] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2298_c2_0b27_cond <= VAR_t16_MUX_uxn_opcodes_h_l2298_c2_0b27_cond;
     t16_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue;
     t16_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output := t16_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2298_c2_0b27] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_500b_uxn_opcodes_h_l2293_l2331_DUPLICATE_50a1 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_500b_uxn_opcodes_h_l2293_l2331_DUPLICATE_50a1_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_500b(
     result,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2298_c2_0b27_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_500b_uxn_opcodes_h_l2293_l2331_DUPLICATE_50a1_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_500b_uxn_opcodes_h_l2293_l2331_DUPLICATE_50a1_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
