-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 2
entity VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_0CLK_4b00ae23 is
port(
 ref_toks_0 : in uint8_t_80;
 var_dim_0 : in unsigned(6 downto 0);
 return_output : out unsigned(7 downto 0));
end VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_0CLK_4b00ae23;
architecture arch of VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_0CLK_4b00ae23 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- uint8_mux128[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570]
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_sel : unsigned(6 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in0 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in1 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in2 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in3 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in4 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in5 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in6 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in7 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in8 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in9 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in10 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in11 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in12 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in13 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in14 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in15 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in16 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in17 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in18 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in19 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in20 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in21 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in22 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in23 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in24 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in25 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in26 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in27 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in28 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in29 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in30 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in31 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in32 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in33 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in34 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in35 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in36 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in37 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in38 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in39 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in40 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in41 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in42 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in43 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in44 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in45 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in46 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in47 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in48 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in49 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in50 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in51 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in52 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in53 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in54 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in55 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in56 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in57 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in58 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in59 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in60 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in61 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in62 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in63 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in64 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in65 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in66 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in67 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in68 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in69 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in70 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in71 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in72 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in73 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in74 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in75 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in76 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in77 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in78 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in79 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in80 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in81 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in82 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in83 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in84 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in85 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in86 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in87 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in88 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in89 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in90 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in91 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in92 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in93 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in94 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in95 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in96 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in97 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in98 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in99 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in100 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in101 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in102 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in103 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in104 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in105 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in106 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in107 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in108 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in109 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in110 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in111 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in112 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in113 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in114 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in115 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in116 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in117 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in118 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in119 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in120 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in121 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in122 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in123 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in124 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in125 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in126 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in127 : unsigned(7 downto 0);
signal uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_return_output : unsigned(7 downto 0);

function uint7_uint7_0( inp : unsigned;
 x : unsigned) return unsigned is

  --variable inp : unsigned(6 downto 0);
  --variable x : unsigned(6 downto 0);
  variable intermediate : unsigned(6 downto 0);
  variable return_output : unsigned(6 downto 0);

begin

    intermediate := (others => '0');
    intermediate(6 downto 0) := unsigned(inp);
    intermediate(6 downto 0) := x;
    
    return_output := intermediate(6 downto 0) ;
    
    return return_output;

end function;


begin

-- SUBMODULE INSTANCES 
-- uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570 : entity work.uint8_mux128_0CLK_9347d63d port map (
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_sel,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in0,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in1,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in2,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in3,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in4,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in5,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in6,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in7,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in8,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in9,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in10,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in11,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in12,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in13,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in14,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in15,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in16,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in17,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in18,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in19,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in20,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in21,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in22,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in23,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in24,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in25,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in26,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in27,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in28,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in29,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in30,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in31,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in32,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in33,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in34,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in35,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in36,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in37,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in38,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in39,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in40,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in41,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in42,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in43,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in44,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in45,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in46,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in47,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in48,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in49,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in50,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in51,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in52,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in53,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in54,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in55,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in56,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in57,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in58,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in59,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in60,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in61,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in62,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in63,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in64,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in65,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in66,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in67,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in68,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in69,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in70,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in71,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in72,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in73,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in74,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in75,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in76,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in77,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in78,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in79,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in80,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in81,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in82,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in83,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in84,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in85,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in86,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in87,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in88,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in89,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in90,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in91,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in92,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in93,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in94,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in95,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in96,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in97,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in98,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in99,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in100,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in101,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in102,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in103,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in104,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in105,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in106,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in107,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in108,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in109,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in110,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in111,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in112,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in113,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in114,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in115,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in116,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in117,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in118,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in119,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in120,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in121,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in122,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in123,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in124,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in125,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in126,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in127,
uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 ref_toks_0,
 var_dim_0,
 -- All submodule outputs
 uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_ref_toks_0 : uint8_t_80;
 variable VAR_var_dim_0 : unsigned(6 downto 0);
 variable VAR_return_output : unsigned(7 downto 0);
 variable VAR_base : uint8_t_80;
 variable VAR_ref_0 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_0_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l14_c10_b745_return_output : unsigned(7 downto 0);
 variable VAR_ref_1 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_1_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l16_c10_eef2_return_output : unsigned(7 downto 0);
 variable VAR_ref_2 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_2_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l18_c10_6767_return_output : unsigned(7 downto 0);
 variable VAR_ref_3 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_3_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l20_c10_a2df_return_output : unsigned(7 downto 0);
 variable VAR_ref_4 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_4_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l22_c10_707a_return_output : unsigned(7 downto 0);
 variable VAR_ref_5 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_5_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l24_c10_16e1_return_output : unsigned(7 downto 0);
 variable VAR_ref_6 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_6_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l26_c10_054d_return_output : unsigned(7 downto 0);
 variable VAR_ref_7 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_7_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l28_c10_880a_return_output : unsigned(7 downto 0);
 variable VAR_ref_8 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_8_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l30_c10_1a13_return_output : unsigned(7 downto 0);
 variable VAR_ref_9 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_9_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l32_c10_99a2_return_output : unsigned(7 downto 0);
 variable VAR_ref_10 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_10_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l34_c11_164f_return_output : unsigned(7 downto 0);
 variable VAR_ref_11 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_11_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l36_c11_b5af_return_output : unsigned(7 downto 0);
 variable VAR_ref_12 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_12_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l38_c11_1b33_return_output : unsigned(7 downto 0);
 variable VAR_ref_13 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_13_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l40_c11_3ac6_return_output : unsigned(7 downto 0);
 variable VAR_ref_14 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_14_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l42_c11_8eaf_return_output : unsigned(7 downto 0);
 variable VAR_ref_15 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_15_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l44_c11_822d_return_output : unsigned(7 downto 0);
 variable VAR_ref_16 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_16_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l46_c11_f3af_return_output : unsigned(7 downto 0);
 variable VAR_ref_17 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_17_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l48_c11_e96c_return_output : unsigned(7 downto 0);
 variable VAR_ref_18 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_18_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l50_c11_260f_return_output : unsigned(7 downto 0);
 variable VAR_ref_19 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_19_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l52_c11_ec9a_return_output : unsigned(7 downto 0);
 variable VAR_ref_20 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_20_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l54_c11_23ed_return_output : unsigned(7 downto 0);
 variable VAR_ref_21 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_21_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l56_c11_0d95_return_output : unsigned(7 downto 0);
 variable VAR_ref_22 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_22_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l58_c11_e496_return_output : unsigned(7 downto 0);
 variable VAR_ref_23 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_23_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l60_c11_242a_return_output : unsigned(7 downto 0);
 variable VAR_ref_24 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_24_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l62_c11_b000_return_output : unsigned(7 downto 0);
 variable VAR_ref_25 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_25_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l64_c11_82a6_return_output : unsigned(7 downto 0);
 variable VAR_ref_26 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_26_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l66_c11_f724_return_output : unsigned(7 downto 0);
 variable VAR_ref_27 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_27_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l68_c11_b484_return_output : unsigned(7 downto 0);
 variable VAR_ref_28 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_28_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l70_c11_8c55_return_output : unsigned(7 downto 0);
 variable VAR_ref_29 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_29_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l72_c11_3735_return_output : unsigned(7 downto 0);
 variable VAR_ref_30 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_30_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l74_c11_8197_return_output : unsigned(7 downto 0);
 variable VAR_ref_31 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_31_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l76_c11_6f4e_return_output : unsigned(7 downto 0);
 variable VAR_ref_32 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_32_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l78_c11_1da0_return_output : unsigned(7 downto 0);
 variable VAR_ref_33 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_33_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l80_c11_855a_return_output : unsigned(7 downto 0);
 variable VAR_ref_34 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_34_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l82_c11_a06e_return_output : unsigned(7 downto 0);
 variable VAR_ref_35 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_35_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l84_c11_fcc4_return_output : unsigned(7 downto 0);
 variable VAR_ref_36 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_36_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l86_c11_a053_return_output : unsigned(7 downto 0);
 variable VAR_ref_37 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_37_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l88_c11_ae5b_return_output : unsigned(7 downto 0);
 variable VAR_ref_38 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_38_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l90_c11_e2d1_return_output : unsigned(7 downto 0);
 variable VAR_ref_39 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_39_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l92_c11_9986_return_output : unsigned(7 downto 0);
 variable VAR_ref_40 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_40_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l94_c11_f7ab_return_output : unsigned(7 downto 0);
 variable VAR_ref_41 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_41_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l96_c11_7e05_return_output : unsigned(7 downto 0);
 variable VAR_ref_42 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_42_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l98_c11_4507_return_output : unsigned(7 downto 0);
 variable VAR_ref_43 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_43_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l100_c11_0472_return_output : unsigned(7 downto 0);
 variable VAR_ref_44 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_44_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l102_c11_f6de_return_output : unsigned(7 downto 0);
 variable VAR_ref_45 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_45_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l104_c11_7bc2_return_output : unsigned(7 downto 0);
 variable VAR_ref_46 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_46_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l106_c11_5d30_return_output : unsigned(7 downto 0);
 variable VAR_ref_47 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_47_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l108_c11_5a1a_return_output : unsigned(7 downto 0);
 variable VAR_ref_48 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_48_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l110_c11_3447_return_output : unsigned(7 downto 0);
 variable VAR_ref_49 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_49_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l112_c11_5ac8_return_output : unsigned(7 downto 0);
 variable VAR_ref_50 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_50_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l114_c11_4a7b_return_output : unsigned(7 downto 0);
 variable VAR_ref_51 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_51_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l116_c11_7ab3_return_output : unsigned(7 downto 0);
 variable VAR_ref_52 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_52_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l118_c11_7d28_return_output : unsigned(7 downto 0);
 variable VAR_ref_53 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_53_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l120_c11_e0a1_return_output : unsigned(7 downto 0);
 variable VAR_ref_54 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_54_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l122_c11_8aa8_return_output : unsigned(7 downto 0);
 variable VAR_ref_55 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_55_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l124_c11_fcd7_return_output : unsigned(7 downto 0);
 variable VAR_ref_56 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_56_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l126_c11_dd80_return_output : unsigned(7 downto 0);
 variable VAR_ref_57 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_57_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l128_c11_2e08_return_output : unsigned(7 downto 0);
 variable VAR_ref_58 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_58_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l130_c11_739f_return_output : unsigned(7 downto 0);
 variable VAR_ref_59 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_59_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l132_c11_01a2_return_output : unsigned(7 downto 0);
 variable VAR_ref_60 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_60_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l134_c11_c28b_return_output : unsigned(7 downto 0);
 variable VAR_ref_61 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_61_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l136_c11_925b_return_output : unsigned(7 downto 0);
 variable VAR_ref_62 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_62_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l138_c11_cb49_return_output : unsigned(7 downto 0);
 variable VAR_ref_63 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_63_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l140_c11_b7d2_return_output : unsigned(7 downto 0);
 variable VAR_ref_64 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_64_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l142_c11_a173_return_output : unsigned(7 downto 0);
 variable VAR_ref_65 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_65_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l144_c11_9329_return_output : unsigned(7 downto 0);
 variable VAR_ref_66 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_66_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l146_c11_e9ff_return_output : unsigned(7 downto 0);
 variable VAR_ref_67 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_67_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l148_c11_aeb1_return_output : unsigned(7 downto 0);
 variable VAR_ref_68 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_68_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l150_c11_e35c_return_output : unsigned(7 downto 0);
 variable VAR_ref_69 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_69_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l152_c11_ce8a_return_output : unsigned(7 downto 0);
 variable VAR_ref_70 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_70_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l154_c11_36ec_return_output : unsigned(7 downto 0);
 variable VAR_ref_71 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_71_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l156_c11_bf2b_return_output : unsigned(7 downto 0);
 variable VAR_ref_72 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_72_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l158_c11_5eeb_return_output : unsigned(7 downto 0);
 variable VAR_ref_73 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_73_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l160_c11_bc2e_return_output : unsigned(7 downto 0);
 variable VAR_ref_74 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_74_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l162_c11_848a_return_output : unsigned(7 downto 0);
 variable VAR_ref_75 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_75_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l164_c11_0f02_return_output : unsigned(7 downto 0);
 variable VAR_ref_76 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_76_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l166_c11_b653_return_output : unsigned(7 downto 0);
 variable VAR_ref_77 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_77_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l168_c11_c1c7_return_output : unsigned(7 downto 0);
 variable VAR_ref_78 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_78_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l170_c11_a033_return_output : unsigned(7 downto 0);
 variable VAR_ref_79 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output : unsigned(7 downto 0);
 variable VAR_sel : unsigned(6 downto 0);
 variable VAR_sel_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l175_c2_ef0f : unsigned(6 downto 0);
 variable VAR_uint7_uint7_0_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l176_c8_dc31_return_output : unsigned(6 downto 0);
 variable VAR_rv : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_sel : unsigned(6 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in0 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in1 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in2 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in3 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in4 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in5 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in6 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in7 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in8 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in9 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in10 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in11 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in12 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in13 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in14 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in15 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in16 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in17 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in18 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in19 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in20 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in21 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in22 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in23 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in24 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in25 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in26 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in27 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in28 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in29 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in30 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in31 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in32 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in33 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in34 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in35 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in36 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in37 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in38 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in39 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in40 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in41 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in42 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in43 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in44 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in45 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in46 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in47 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in48 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in49 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in50 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in51 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in52 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in53 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in54 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in55 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in56 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in57 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in58 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in59 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in60 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in61 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in62 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in63 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in64 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in65 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in66 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in67 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in68 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in69 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in70 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in71 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in72 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in73 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in74 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in75 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in76 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in77 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in78 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in79 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in80 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in81 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in82 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in83 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in84 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in85 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in86 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in87 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in88 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in89 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in90 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in91 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in92 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in93 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in94 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in95 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in96 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in97 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in98 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in99 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in100 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in101 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in102 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in103 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in104 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in105 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in106 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in107 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in108 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in109 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in110 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in111 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in112 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in113 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in114 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in115 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in116 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in117 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in118 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in119 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in120 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in121 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in122 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in123 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in124 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in125 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in126 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in127 : unsigned(7 downto 0);
 variable VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_return_output : unsigned(7 downto 0);
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sel_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l175_c2_ef0f := resize(to_unsigned(0, 1), 7);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_ref_toks_0 := ref_toks_0;
     VAR_var_dim_0 := var_dim_0;

     -- Submodule level 0
     -- CONST_REF_RD_uint8_t_uint8_t_80_9_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l32_c10_99a2] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_9_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l32_c10_99a2_return_output := VAR_ref_toks_0(9);

     -- CONST_REF_RD_uint8_t_uint8_t_80_28_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l70_c11_8c55] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_28_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l70_c11_8c55_return_output := VAR_ref_toks_0(28);

     -- CONST_REF_RD_uint8_t_uint8_t_80_53_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l120_c11_e0a1] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_53_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l120_c11_e0a1_return_output := VAR_ref_toks_0(53);

     -- CONST_REF_RD_uint8_t_uint8_t_80_5_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l24_c10_16e1] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_5_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l24_c10_16e1_return_output := VAR_ref_toks_0(5);

     -- CONST_REF_RD_uint8_t_uint8_t_80_76_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l166_c11_b653] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_76_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l166_c11_b653_return_output := VAR_ref_toks_0(76);

     -- CONST_REF_RD_uint8_t_uint8_t_80_10_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l34_c11_164f] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_10_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l34_c11_164f_return_output := VAR_ref_toks_0(10);

     -- CONST_REF_RD_uint8_t_uint8_t_80_32_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l78_c11_1da0] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_32_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l78_c11_1da0_return_output := VAR_ref_toks_0(32);

     -- CONST_REF_RD_uint8_t_uint8_t_80_45_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l104_c11_7bc2] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_45_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l104_c11_7bc2_return_output := VAR_ref_toks_0(45);

     -- CONST_REF_RD_uint8_t_uint8_t_80_39_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l92_c11_9986] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_39_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l92_c11_9986_return_output := VAR_ref_toks_0(39);

     -- CONST_REF_RD_uint8_t_uint8_t_80_65_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l144_c11_9329] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_65_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l144_c11_9329_return_output := VAR_ref_toks_0(65);

     -- CONST_REF_RD_uint8_t_uint8_t_80_62_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l138_c11_cb49] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_62_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l138_c11_cb49_return_output := VAR_ref_toks_0(62);

     -- CONST_REF_RD_uint8_t_uint8_t_80_34_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l82_c11_a06e] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_34_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l82_c11_a06e_return_output := VAR_ref_toks_0(34);

     -- CONST_REF_RD_uint8_t_uint8_t_80_18_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l50_c11_260f] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_18_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l50_c11_260f_return_output := VAR_ref_toks_0(18);

     -- CONST_REF_RD_uint8_t_uint8_t_80_13_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l40_c11_3ac6] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_13_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l40_c11_3ac6_return_output := VAR_ref_toks_0(13);

     -- CONST_REF_RD_uint8_t_uint8_t_80_3_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l20_c10_a2df] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_3_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l20_c10_a2df_return_output := VAR_ref_toks_0(3);

     -- CONST_REF_RD_uint8_t_uint8_t_80_55_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l124_c11_fcd7] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_55_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l124_c11_fcd7_return_output := VAR_ref_toks_0(55);

     -- CONST_REF_RD_uint8_t_uint8_t_80_0_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l14_c10_b745] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_0_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l14_c10_b745_return_output := VAR_ref_toks_0(0);

     -- CONST_REF_RD_uint8_t_uint8_t_80_22_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l58_c11_e496] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_22_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l58_c11_e496_return_output := VAR_ref_toks_0(22);

     -- CONST_REF_RD_uint8_t_uint8_t_80_21_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l56_c11_0d95] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_21_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l56_c11_0d95_return_output := VAR_ref_toks_0(21);

     -- CONST_REF_RD_uint8_t_uint8_t_80_26_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l66_c11_f724] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_26_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l66_c11_f724_return_output := VAR_ref_toks_0(26);

     -- CONST_REF_RD_uint8_t_uint8_t_80_69_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l152_c11_ce8a] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_69_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l152_c11_ce8a_return_output := VAR_ref_toks_0(69);

     -- CONST_REF_RD_uint8_t_uint8_t_80_74_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l162_c11_848a] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_74_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l162_c11_848a_return_output := VAR_ref_toks_0(74);

     -- CONST_REF_RD_uint8_t_uint8_t_80_31_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l76_c11_6f4e] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_31_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l76_c11_6f4e_return_output := VAR_ref_toks_0(31);

     -- CONST_REF_RD_uint8_t_uint8_t_80_68_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l150_c11_e35c] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_68_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l150_c11_e35c_return_output := VAR_ref_toks_0(68);

     -- CONST_REF_RD_uint8_t_uint8_t_80_37_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l88_c11_ae5b] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_37_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l88_c11_ae5b_return_output := VAR_ref_toks_0(37);

     -- CONST_REF_RD_uint8_t_uint8_t_80_49_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l112_c11_5ac8] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_49_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l112_c11_5ac8_return_output := VAR_ref_toks_0(49);

     -- CONST_REF_RD_uint8_t_uint8_t_80_60_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l134_c11_c28b] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_60_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l134_c11_c28b_return_output := VAR_ref_toks_0(60);

     -- CONST_REF_RD_uint8_t_uint8_t_80_73_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l160_c11_bc2e] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_73_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l160_c11_bc2e_return_output := VAR_ref_toks_0(73);

     -- CONST_REF_RD_uint8_t_uint8_t_80_54_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l122_c11_8aa8] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_54_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l122_c11_8aa8_return_output := VAR_ref_toks_0(54);

     -- CONST_REF_RD_uint8_t_uint8_t_80_61_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l136_c11_925b] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_61_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l136_c11_925b_return_output := VAR_ref_toks_0(61);

     -- CONST_REF_RD_uint8_t_uint8_t_80_64_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l142_c11_a173] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_64_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l142_c11_a173_return_output := VAR_ref_toks_0(64);

     -- CONST_REF_RD_uint8_t_uint8_t_80_41_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l96_c11_7e05] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_41_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l96_c11_7e05_return_output := VAR_ref_toks_0(41);

     -- CONST_REF_RD_uint8_t_uint8_t_80_63_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l140_c11_b7d2] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_63_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l140_c11_b7d2_return_output := VAR_ref_toks_0(63);

     -- CONST_REF_RD_uint8_t_uint8_t_80_56_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l126_c11_dd80] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_56_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l126_c11_dd80_return_output := VAR_ref_toks_0(56);

     -- CONST_REF_RD_uint8_t_uint8_t_80_2_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l18_c10_6767] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_2_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l18_c10_6767_return_output := VAR_ref_toks_0(2);

     -- CONST_REF_RD_uint8_t_uint8_t_80_77_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l168_c11_c1c7] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_77_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l168_c11_c1c7_return_output := VAR_ref_toks_0(77);

     -- CONST_REF_RD_uint8_t_uint8_t_80_1_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l16_c10_eef2] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_1_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l16_c10_eef2_return_output := VAR_ref_toks_0(1);

     -- CONST_REF_RD_uint8_t_uint8_t_80_8_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l30_c10_1a13] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_8_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l30_c10_1a13_return_output := VAR_ref_toks_0(8);

     -- CONST_REF_RD_uint8_t_uint8_t_80_58_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l130_c11_739f] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_58_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l130_c11_739f_return_output := VAR_ref_toks_0(58);

     -- CONST_REF_RD_uint8_t_uint8_t_80_75_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l164_c11_0f02] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_75_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l164_c11_0f02_return_output := VAR_ref_toks_0(75);

     -- CONST_REF_RD_uint8_t_uint8_t_80_57_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l128_c11_2e08] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_57_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l128_c11_2e08_return_output := VAR_ref_toks_0(57);

     -- CONST_REF_RD_uint8_t_uint8_t_80_70_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l154_c11_36ec] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_70_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l154_c11_36ec_return_output := VAR_ref_toks_0(70);

     -- CONST_REF_RD_uint8_t_uint8_t_80_29_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l72_c11_3735] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_29_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l72_c11_3735_return_output := VAR_ref_toks_0(29);

     -- CONST_REF_RD_uint8_t_uint8_t_80_14_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l42_c11_8eaf] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_14_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l42_c11_8eaf_return_output := VAR_ref_toks_0(14);

     -- CONST_REF_RD_uint8_t_uint8_t_80_46_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l106_c11_5d30] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_46_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l106_c11_5d30_return_output := VAR_ref_toks_0(46);

     -- CONST_REF_RD_uint8_t_uint8_t_80_16_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l46_c11_f3af] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_16_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l46_c11_f3af_return_output := VAR_ref_toks_0(16);

     -- CONST_REF_RD_uint8_t_uint8_t_80_24_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l62_c11_b000] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_24_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l62_c11_b000_return_output := VAR_ref_toks_0(24);

     -- CONST_REF_RD_uint8_t_uint8_t_80_40_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l94_c11_f7ab] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_40_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l94_c11_f7ab_return_output := VAR_ref_toks_0(40);

     -- CONST_REF_RD_uint8_t_uint8_t_80_72_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l158_c11_5eeb] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_72_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l158_c11_5eeb_return_output := VAR_ref_toks_0(72);

     -- CONST_REF_RD_uint8_t_uint8_t_80_27_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l68_c11_b484] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_27_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l68_c11_b484_return_output := VAR_ref_toks_0(27);

     -- CONST_REF_RD_uint8_t_uint8_t_80_66_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l146_c11_e9ff] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_66_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l146_c11_e9ff_return_output := VAR_ref_toks_0(66);

     -- CONST_REF_RD_uint8_t_uint8_t_80_47_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l108_c11_5a1a] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_47_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l108_c11_5a1a_return_output := VAR_ref_toks_0(47);

     -- CONST_REF_RD_uint8_t_uint8_t_80_33_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l80_c11_855a] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_33_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l80_c11_855a_return_output := VAR_ref_toks_0(33);

     -- CONST_REF_RD_uint8_t_uint8_t_80_48_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l110_c11_3447] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_48_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l110_c11_3447_return_output := VAR_ref_toks_0(48);

     -- CONST_REF_RD_uint8_t_uint8_t_80_17_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l48_c11_e96c] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_17_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l48_c11_e96c_return_output := VAR_ref_toks_0(17);

     -- CONST_REF_RD_uint8_t_uint8_t_80_25_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l64_c11_82a6] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_25_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l64_c11_82a6_return_output := VAR_ref_toks_0(25);

     -- CONST_REF_RD_uint8_t_uint8_t_80_6_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l26_c10_054d] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_6_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l26_c10_054d_return_output := VAR_ref_toks_0(6);

     -- CONST_REF_RD_uint8_t_uint8_t_80_23_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l60_c11_242a] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_23_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l60_c11_242a_return_output := VAR_ref_toks_0(23);

     -- CONST_REF_RD_uint8_t_uint8_t_80_67_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l148_c11_aeb1] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_67_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l148_c11_aeb1_return_output := VAR_ref_toks_0(67);

     -- CONST_REF_RD_uint8_t_uint8_t_80_78_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l170_c11_a033] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_78_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l170_c11_a033_return_output := VAR_ref_toks_0(78);

     -- CONST_REF_RD_uint8_t_uint8_t_80_79_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output := VAR_ref_toks_0(79);

     -- CONST_REF_RD_uint8_t_uint8_t_80_43_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l100_c11_0472] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_43_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l100_c11_0472_return_output := VAR_ref_toks_0(43);

     -- CONST_REF_RD_uint8_t_uint8_t_80_59_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l132_c11_01a2] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_59_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l132_c11_01a2_return_output := VAR_ref_toks_0(59);

     -- CONST_REF_RD_uint8_t_uint8_t_80_4_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l22_c10_707a] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_4_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l22_c10_707a_return_output := VAR_ref_toks_0(4);

     -- CONST_REF_RD_uint8_t_uint8_t_80_50_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l114_c11_4a7b] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_50_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l114_c11_4a7b_return_output := VAR_ref_toks_0(50);

     -- uint7_uint7_0[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l176_c8_dc31] LATENCY=0
     VAR_uint7_uint7_0_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l176_c8_dc31_return_output := uint7_uint7_0(
     VAR_sel_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l175_c2_ef0f,
     VAR_var_dim_0);

     -- CONST_REF_RD_uint8_t_uint8_t_80_19_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l52_c11_ec9a] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_19_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l52_c11_ec9a_return_output := VAR_ref_toks_0(19);

     -- CONST_REF_RD_uint8_t_uint8_t_80_71_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l156_c11_bf2b] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_71_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l156_c11_bf2b_return_output := VAR_ref_toks_0(71);

     -- CONST_REF_RD_uint8_t_uint8_t_80_12_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l38_c11_1b33] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_12_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l38_c11_1b33_return_output := VAR_ref_toks_0(12);

     -- CONST_REF_RD_uint8_t_uint8_t_80_15_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l44_c11_822d] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_15_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l44_c11_822d_return_output := VAR_ref_toks_0(15);

     -- CONST_REF_RD_uint8_t_uint8_t_80_42_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l98_c11_4507] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_42_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l98_c11_4507_return_output := VAR_ref_toks_0(42);

     -- CONST_REF_RD_uint8_t_uint8_t_80_20_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l54_c11_23ed] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_20_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l54_c11_23ed_return_output := VAR_ref_toks_0(20);

     -- CONST_REF_RD_uint8_t_uint8_t_80_30_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l74_c11_8197] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_30_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l74_c11_8197_return_output := VAR_ref_toks_0(30);

     -- CONST_REF_RD_uint8_t_uint8_t_80_52_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l118_c11_7d28] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_52_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l118_c11_7d28_return_output := VAR_ref_toks_0(52);

     -- CONST_REF_RD_uint8_t_uint8_t_80_36_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l86_c11_a053] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_36_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l86_c11_a053_return_output := VAR_ref_toks_0(36);

     -- CONST_REF_RD_uint8_t_uint8_t_80_35_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l84_c11_fcc4] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_35_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l84_c11_fcc4_return_output := VAR_ref_toks_0(35);

     -- CONST_REF_RD_uint8_t_uint8_t_80_7_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l28_c10_880a] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_7_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l28_c10_880a_return_output := VAR_ref_toks_0(7);

     -- CONST_REF_RD_uint8_t_uint8_t_80_11_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l36_c11_b5af] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_11_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l36_c11_b5af_return_output := VAR_ref_toks_0(11);

     -- CONST_REF_RD_uint8_t_uint8_t_80_51_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l116_c11_7ab3] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_51_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l116_c11_7ab3_return_output := VAR_ref_toks_0(51);

     -- CONST_REF_RD_uint8_t_uint8_t_80_38_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l90_c11_e2d1] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_38_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l90_c11_e2d1_return_output := VAR_ref_toks_0(38);

     -- CONST_REF_RD_uint8_t_uint8_t_80_44_d41d[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l102_c11_f6de] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_80_44_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l102_c11_f6de_return_output := VAR_ref_toks_0(44);

     -- Submodule level 1
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in0 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_0_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l14_c10_b745_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in10 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_10_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l34_c11_164f_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in11 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_11_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l36_c11_b5af_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in12 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_12_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l38_c11_1b33_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in13 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_13_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l40_c11_3ac6_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in14 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_14_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l42_c11_8eaf_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in15 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_15_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l44_c11_822d_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in16 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_16_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l46_c11_f3af_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in17 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_17_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l48_c11_e96c_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in18 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_18_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l50_c11_260f_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in19 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_19_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l52_c11_ec9a_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in1 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_1_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l16_c10_eef2_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in20 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_20_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l54_c11_23ed_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in21 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_21_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l56_c11_0d95_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in22 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_22_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l58_c11_e496_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in23 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_23_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l60_c11_242a_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in24 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_24_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l62_c11_b000_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in25 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_25_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l64_c11_82a6_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in26 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_26_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l66_c11_f724_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in27 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_27_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l68_c11_b484_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in28 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_28_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l70_c11_8c55_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in29 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_29_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l72_c11_3735_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in2 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_2_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l18_c10_6767_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in30 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_30_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l74_c11_8197_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in31 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_31_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l76_c11_6f4e_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in32 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_32_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l78_c11_1da0_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in33 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_33_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l80_c11_855a_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in34 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_34_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l82_c11_a06e_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in35 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_35_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l84_c11_fcc4_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in36 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_36_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l86_c11_a053_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in37 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_37_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l88_c11_ae5b_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in38 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_38_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l90_c11_e2d1_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in39 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_39_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l92_c11_9986_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in3 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_3_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l20_c10_a2df_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in40 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_40_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l94_c11_f7ab_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in41 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_41_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l96_c11_7e05_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in42 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_42_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l98_c11_4507_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in43 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_43_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l100_c11_0472_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in44 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_44_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l102_c11_f6de_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in45 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_45_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l104_c11_7bc2_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in46 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_46_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l106_c11_5d30_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in47 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_47_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l108_c11_5a1a_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in48 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_48_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l110_c11_3447_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in49 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_49_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l112_c11_5ac8_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in4 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_4_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l22_c10_707a_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in50 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_50_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l114_c11_4a7b_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in51 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_51_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l116_c11_7ab3_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in52 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_52_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l118_c11_7d28_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in53 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_53_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l120_c11_e0a1_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in54 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_54_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l122_c11_8aa8_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in55 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_55_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l124_c11_fcd7_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in56 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_56_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l126_c11_dd80_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in57 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_57_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l128_c11_2e08_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in58 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_58_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l130_c11_739f_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in59 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_59_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l132_c11_01a2_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in5 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_5_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l24_c10_16e1_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in60 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_60_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l134_c11_c28b_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in61 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_61_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l136_c11_925b_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in62 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_62_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l138_c11_cb49_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in63 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_63_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l140_c11_b7d2_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in64 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_64_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l142_c11_a173_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in65 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_65_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l144_c11_9329_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in66 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_66_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l146_c11_e9ff_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in67 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_67_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l148_c11_aeb1_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in68 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_68_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l150_c11_e35c_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in69 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_69_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l152_c11_ce8a_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in6 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_6_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l26_c10_054d_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in70 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_70_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l154_c11_36ec_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in71 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_71_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l156_c11_bf2b_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in72 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_72_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l158_c11_5eeb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in73 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_73_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l160_c11_bc2e_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in74 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_74_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l162_c11_848a_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in75 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_75_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l164_c11_0f02_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in76 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_76_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l166_c11_b653_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in77 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_77_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l168_c11_c1c7_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in78 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_78_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l170_c11_a033_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in100 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in101 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in102 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in103 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in104 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in105 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in106 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in107 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in108 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in109 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in110 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in111 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in112 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in113 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in114 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in115 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in116 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in117 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in118 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in119 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in120 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in121 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in122 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in123 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in124 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in125 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in126 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in127 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in79 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in80 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in81 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in82 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in83 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in84 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in85 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in86 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in87 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in88 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in89 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in90 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in91 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in92 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in93 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in94 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in95 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in96 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in97 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in98 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in99 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_79_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l172_c11_2feb_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in7 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_7_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l28_c10_880a_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in8 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_8_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l30_c10_1a13_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in9 := VAR_CONST_REF_RD_uint8_t_uint8_t_80_9_d41d_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l32_c10_99a2_return_output;
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_sel := VAR_uint7_uint7_0_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l176_c8_dc31_return_output;
     -- uint8_mux128[VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570] LATENCY=0
     -- Inputs
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_sel <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_sel;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in0 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in0;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in1 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in1;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in2 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in2;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in3 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in3;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in4 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in4;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in5 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in5;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in6 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in6;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in7 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in7;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in8 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in8;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in9 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in9;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in10 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in10;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in11 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in11;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in12 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in12;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in13 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in13;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in14 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in14;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in15 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in15;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in16 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in16;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in17 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in17;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in18 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in18;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in19 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in19;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in20 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in20;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in21 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in21;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in22 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in22;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in23 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in23;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in24 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in24;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in25 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in25;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in26 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in26;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in27 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in27;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in28 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in28;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in29 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in29;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in30 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in30;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in31 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in31;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in32 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in32;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in33 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in33;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in34 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in34;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in35 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in35;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in36 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in36;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in37 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in37;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in38 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in38;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in39 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in39;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in40 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in40;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in41 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in41;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in42 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in42;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in43 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in43;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in44 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in44;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in45 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in45;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in46 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in46;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in47 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in47;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in48 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in48;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in49 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in49;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in50 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in50;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in51 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in51;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in52 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in52;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in53 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in53;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in54 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in54;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in55 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in55;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in56 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in56;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in57 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in57;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in58 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in58;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in59 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in59;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in60 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in60;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in61 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in61;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in62 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in62;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in63 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in63;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in64 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in64;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in65 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in65;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in66 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in66;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in67 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in67;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in68 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in68;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in69 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in69;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in70 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in70;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in71 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in71;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in72 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in72;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in73 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in73;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in74 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in74;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in75 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in75;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in76 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in76;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in77 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in77;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in78 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in78;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in79 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in79;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in80 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in80;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in81 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in81;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in82 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in82;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in83 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in83;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in84 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in84;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in85 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in85;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in86 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in86;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in87 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in87;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in88 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in88;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in89 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in89;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in90 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in90;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in91 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in91;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in92 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in92;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in93 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in93;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in94 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in94;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in95 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in95;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in96 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in96;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in97 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in97;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in98 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in98;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in99 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in99;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in100 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in100;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in101 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in101;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in102 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in102;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in103 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in103;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in104 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in104;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in105 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in105;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in106 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in106;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in107 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in107;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in108 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in108;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in109 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in109;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in110 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in110;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in111 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in111;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in112 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in112;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in113 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in113;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in114 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in114;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in115 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in115;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in116 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in116;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in117 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in117;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in118 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in118;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in119 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in119;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in120 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in120;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in121 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in121;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in122 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in122;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in123 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in123;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in124 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in124;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in125 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in125;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in126 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in126;
     uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in127 <= VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_in127;
     -- Outputs
     VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_return_output := uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_return_output;

     -- Submodule level 2
     VAR_return_output := VAR_uint8_mux128_VAR_REF_RD_uint8_t_uint8_t_80_VAR_d41d_c_l179_c7_4570_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
