-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity lth_0CLK_85d5529e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end lth_0CLK_85d5529e;
architecture arch of lth_0CLK_85d5529e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1800_c6_0818]
signal BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1800_c1_07d6]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1800_c2_414f]
signal n8_MUX_uxn_opcodes_h_l1800_c2_414f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1800_c2_414f_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1800_c2_414f]
signal t8_MUX_uxn_opcodes_h_l1800_c2_414f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1800_c2_414f_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1800_c2_414f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1800_c2_414f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1800_c2_414f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1800_c2_414f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1800_c2_414f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1800_c2_414f]
signal result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1801_c3_b0c0[uxn_opcodes_h_l1801_c3_b0c0]
signal printf_uxn_opcodes_h_l1801_c3_b0c0_uxn_opcodes_h_l1801_c3_b0c0_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1805_c11_7fed]
signal BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1805_c7_517b]
signal n8_MUX_uxn_opcodes_h_l1805_c7_517b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1805_c7_517b_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1805_c7_517b]
signal t8_MUX_uxn_opcodes_h_l1805_c7_517b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1805_c7_517b_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1805_c7_517b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1805_c7_517b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1805_c7_517b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1805_c7_517b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1805_c7_517b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1805_c7_517b]
signal result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1808_c11_3ff5]
signal BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1808_c7_e477]
signal n8_MUX_uxn_opcodes_h_l1808_c7_e477_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1808_c7_e477_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1808_c7_e477]
signal t8_MUX_uxn_opcodes_h_l1808_c7_e477_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1808_c7_e477_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1808_c7_e477]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1808_c7_e477]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1808_c7_e477]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1808_c7_e477]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1808_c7_e477]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1808_c7_e477]
signal result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1811_c11_63ae]
signal BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1811_c7_760f]
signal n8_MUX_uxn_opcodes_h_l1811_c7_760f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1811_c7_760f_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1811_c7_760f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1811_c7_760f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1811_c7_760f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1811_c7_760f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1811_c7_760f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1811_c7_760f]
signal result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1814_c30_a6ce]
signal sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_return_output : signed(3 downto 0);

-- BIN_OP_LT[uxn_opcodes_h_l1817_c21_c087]
signal BIN_OP_LT_uxn_opcodes_h_l1817_c21_c087_left : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l1817_c21_c087_right : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l1817_c21_c087_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1817_c21_6dee]
signal MUX_uxn_opcodes_h_l1817_c21_6dee_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1817_c21_6dee_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1817_c21_6dee_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1817_c21_6dee_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1819_c11_206f]
signal BIN_OP_EQ_uxn_opcodes_h_l1819_c11_206f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1819_c11_206f_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1819_c11_206f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1819_c7_7e65]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1819_c7_7e65]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1819_c7_7e65]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_4e73( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818
BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_left,
BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_right,
BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_return_output);

-- n8_MUX_uxn_opcodes_h_l1800_c2_414f
n8_MUX_uxn_opcodes_h_l1800_c2_414f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1800_c2_414f_cond,
n8_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue,
n8_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse,
n8_MUX_uxn_opcodes_h_l1800_c2_414f_return_output);

-- t8_MUX_uxn_opcodes_h_l1800_c2_414f
t8_MUX_uxn_opcodes_h_l1800_c2_414f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1800_c2_414f_cond,
t8_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue,
t8_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse,
t8_MUX_uxn_opcodes_h_l1800_c2_414f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f
result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f
result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f
result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f
result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_return_output);

-- printf_uxn_opcodes_h_l1801_c3_b0c0_uxn_opcodes_h_l1801_c3_b0c0
printf_uxn_opcodes_h_l1801_c3_b0c0_uxn_opcodes_h_l1801_c3_b0c0 : entity work.printf_uxn_opcodes_h_l1801_c3_b0c0_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1801_c3_b0c0_uxn_opcodes_h_l1801_c3_b0c0_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed
BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_left,
BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_right,
BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_return_output);

-- n8_MUX_uxn_opcodes_h_l1805_c7_517b
n8_MUX_uxn_opcodes_h_l1805_c7_517b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1805_c7_517b_cond,
n8_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue,
n8_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse,
n8_MUX_uxn_opcodes_h_l1805_c7_517b_return_output);

-- t8_MUX_uxn_opcodes_h_l1805_c7_517b
t8_MUX_uxn_opcodes_h_l1805_c7_517b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1805_c7_517b_cond,
t8_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue,
t8_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse,
t8_MUX_uxn_opcodes_h_l1805_c7_517b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b
result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b
result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b
result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b
result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5
BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_left,
BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_right,
BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_return_output);

-- n8_MUX_uxn_opcodes_h_l1808_c7_e477
n8_MUX_uxn_opcodes_h_l1808_c7_e477 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1808_c7_e477_cond,
n8_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue,
n8_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse,
n8_MUX_uxn_opcodes_h_l1808_c7_e477_return_output);

-- t8_MUX_uxn_opcodes_h_l1808_c7_e477
t8_MUX_uxn_opcodes_h_l1808_c7_e477 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1808_c7_e477_cond,
t8_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue,
t8_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse,
t8_MUX_uxn_opcodes_h_l1808_c7_e477_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477
result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477
result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477
result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477
result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477
result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_cond,
result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae
BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_left,
BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_right,
BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_return_output);

-- n8_MUX_uxn_opcodes_h_l1811_c7_760f
n8_MUX_uxn_opcodes_h_l1811_c7_760f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1811_c7_760f_cond,
n8_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue,
n8_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse,
n8_MUX_uxn_opcodes_h_l1811_c7_760f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f
result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f
result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f
result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f
result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce
sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_ins,
sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_x,
sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_y,
sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_return_output);

-- BIN_OP_LT_uxn_opcodes_h_l1817_c21_c087
BIN_OP_LT_uxn_opcodes_h_l1817_c21_c087 : entity work.BIN_OP_LT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_LT_uxn_opcodes_h_l1817_c21_c087_left,
BIN_OP_LT_uxn_opcodes_h_l1817_c21_c087_right,
BIN_OP_LT_uxn_opcodes_h_l1817_c21_c087_return_output);

-- MUX_uxn_opcodes_h_l1817_c21_6dee
MUX_uxn_opcodes_h_l1817_c21_6dee : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1817_c21_6dee_cond,
MUX_uxn_opcodes_h_l1817_c21_6dee_iftrue,
MUX_uxn_opcodes_h_l1817_c21_6dee_iffalse,
MUX_uxn_opcodes_h_l1817_c21_6dee_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1819_c11_206f
BIN_OP_EQ_uxn_opcodes_h_l1819_c11_206f : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1819_c11_206f_left,
BIN_OP_EQ_uxn_opcodes_h_l1819_c11_206f_right,
BIN_OP_EQ_uxn_opcodes_h_l1819_c11_206f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65
result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65
result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65
result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_return_output,
 n8_MUX_uxn_opcodes_h_l1800_c2_414f_return_output,
 t8_MUX_uxn_opcodes_h_l1800_c2_414f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_return_output,
 n8_MUX_uxn_opcodes_h_l1805_c7_517b_return_output,
 t8_MUX_uxn_opcodes_h_l1805_c7_517b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_return_output,
 n8_MUX_uxn_opcodes_h_l1808_c7_e477_return_output,
 t8_MUX_uxn_opcodes_h_l1808_c7_e477_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_return_output,
 n8_MUX_uxn_opcodes_h_l1811_c7_760f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_return_output,
 sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_return_output,
 BIN_OP_LT_uxn_opcodes_h_l1817_c21_c087_return_output,
 MUX_uxn_opcodes_h_l1817_c21_6dee_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1819_c11_206f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1805_c7_517b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1800_c2_414f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1800_c2_414f_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1805_c7_517b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1800_c2_414f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1800_c2_414f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1802_c3_bb62 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1801_c3_b0c0_uxn_opcodes_h_l1801_c3_b0c0_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1808_c7_e477_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1805_c7_517b_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1808_c7_e477_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1805_c7_517b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1806_c3_e252 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1811_c7_760f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1808_c7_e477_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1808_c7_e477_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1811_c7_760f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1816_c3_3d36 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1817_c21_6dee_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1817_c21_6dee_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1817_c21_6dee_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_c087_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_c087_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_c087_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1817_c21_6dee_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_206f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_206f_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_206f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1808_l1800_l1805_l1819_DUPLICATE_0b55_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1808_l1800_l1805_l1819_DUPLICATE_4978_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1808_l1800_l1811_l1805_DUPLICATE_e839_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1808_l1800_l1811_l1805_DUPLICATE_cf9d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1808_l1811_l1805_l1819_DUPLICATE_dbfa_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1808_l1811_DUPLICATE_672a_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l1796_l1825_DUPLICATE_b86c_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1817_c21_6dee_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_iffalse := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1817_c21_6dee_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_206f_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1802_c3_bb62 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1802_c3_bb62;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1816_c3_3d36 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1816_c3_3d36;
     VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1806_c3_e252 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1806_c3_e252;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_right := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_206f_left := VAR_phase;
     VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_c087_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_c087_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse := t8;
     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1808_l1811_DUPLICATE_672a LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1808_l1811_DUPLICATE_672a_return_output := result.stack_address_sp_offset;

     -- BIN_OP_LT[uxn_opcodes_h_l1817_c21_c087] LATENCY=0
     -- Inputs
     BIN_OP_LT_uxn_opcodes_h_l1817_c21_c087_left <= VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_c087_left;
     BIN_OP_LT_uxn_opcodes_h_l1817_c21_c087_right <= VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_c087_right;
     -- Outputs
     VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_c087_return_output := BIN_OP_LT_uxn_opcodes_h_l1817_c21_c087_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1808_l1811_l1805_l1819_DUPLICATE_dbfa LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1808_l1811_l1805_l1819_DUPLICATE_dbfa_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1808_l1800_l1805_l1819_DUPLICATE_0b55 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1808_l1800_l1805_l1819_DUPLICATE_0b55_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1800_c6_0818] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_left;
     BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_return_output := BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1808_c11_3ff5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_left;
     BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_return_output := BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1811_c11_63ae] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_left;
     BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_return_output := BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1808_l1800_l1811_l1805_DUPLICATE_e839 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1808_l1800_l1811_l1805_DUPLICATE_e839_return_output := result.sp_relative_shift;

     -- sp_relative_shift[uxn_opcodes_h_l1814_c30_a6ce] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_ins;
     sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_x;
     sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_return_output := sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1805_c11_7fed] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_left;
     BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_return_output := BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1819_c11_206f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1819_c11_206f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_206f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1819_c11_206f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_206f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_206f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1819_c11_206f_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1808_l1800_l1805_l1819_DUPLICATE_4978 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1808_l1800_l1805_l1819_DUPLICATE_4978_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1808_l1800_l1811_l1805_DUPLICATE_cf9d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1808_l1800_l1811_l1805_DUPLICATE_cf9d_return_output := result.u8_value;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1800_c2_414f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1800_c2_414f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_0818_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1805_c7_517b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1805_c7_517b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_7fed_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1808_c7_e477_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1808_c7_e477_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_3ff5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1811_c7_760f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_63ae_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_206f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_206f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_206f_return_output;
     VAR_MUX_uxn_opcodes_h_l1817_c21_6dee_cond := VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_c087_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1808_l1800_l1811_l1805_DUPLICATE_e839_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1808_l1800_l1811_l1805_DUPLICATE_e839_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1808_l1800_l1811_l1805_DUPLICATE_e839_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1808_l1800_l1811_l1805_DUPLICATE_e839_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1808_l1811_l1805_l1819_DUPLICATE_dbfa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1808_l1811_l1805_l1819_DUPLICATE_dbfa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1808_l1811_l1805_l1819_DUPLICATE_dbfa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1808_l1811_l1805_l1819_DUPLICATE_dbfa_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1808_l1800_l1805_l1819_DUPLICATE_4978_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1808_l1800_l1805_l1819_DUPLICATE_4978_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1808_l1800_l1805_l1819_DUPLICATE_4978_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1808_l1800_l1805_l1819_DUPLICATE_4978_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1808_l1800_l1805_l1819_DUPLICATE_0b55_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1808_l1800_l1805_l1819_DUPLICATE_0b55_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1808_l1800_l1805_l1819_DUPLICATE_0b55_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1808_l1800_l1805_l1819_DUPLICATE_0b55_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1808_l1811_DUPLICATE_672a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1808_l1811_DUPLICATE_672a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1808_l1800_l1811_l1805_DUPLICATE_cf9d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1808_l1800_l1811_l1805_DUPLICATE_cf9d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1808_l1800_l1811_l1805_DUPLICATE_cf9d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1808_l1800_l1811_l1805_DUPLICATE_cf9d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_a6ce_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1819_c7_7e65] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1811_c7_760f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_return_output;

     -- t8_MUX[uxn_opcodes_h_l1808_c7_e477] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1808_c7_e477_cond <= VAR_t8_MUX_uxn_opcodes_h_l1808_c7_e477_cond;
     t8_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue;
     t8_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1808_c7_e477_return_output := t8_MUX_uxn_opcodes_h_l1808_c7_e477_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1800_c1_07d6] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1819_c7_7e65] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_return_output;

     -- n8_MUX[uxn_opcodes_h_l1811_c7_760f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1811_c7_760f_cond <= VAR_n8_MUX_uxn_opcodes_h_l1811_c7_760f_cond;
     n8_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue;
     n8_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1811_c7_760f_return_output := n8_MUX_uxn_opcodes_h_l1811_c7_760f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1819_c7_7e65] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_return_output;

     -- MUX[uxn_opcodes_h_l1817_c21_6dee] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1817_c21_6dee_cond <= VAR_MUX_uxn_opcodes_h_l1817_c21_6dee_cond;
     MUX_uxn_opcodes_h_l1817_c21_6dee_iftrue <= VAR_MUX_uxn_opcodes_h_l1817_c21_6dee_iftrue;
     MUX_uxn_opcodes_h_l1817_c21_6dee_iffalse <= VAR_MUX_uxn_opcodes_h_l1817_c21_6dee_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1817_c21_6dee_return_output := MUX_uxn_opcodes_h_l1817_c21_6dee_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1811_c7_760f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue := VAR_MUX_uxn_opcodes_h_l1817_c21_6dee_return_output;
     VAR_printf_uxn_opcodes_h_l1801_c3_b0c0_uxn_opcodes_h_l1801_c3_b0c0_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_07d6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1811_c7_760f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_7e65_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_7e65_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_7e65_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_760f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_760f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1808_c7_e477_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1808_c7_e477] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1811_c7_760f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1811_c7_760f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_return_output;

     -- printf_uxn_opcodes_h_l1801_c3_b0c0[uxn_opcodes_h_l1801_c3_b0c0] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1801_c3_b0c0_uxn_opcodes_h_l1801_c3_b0c0_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1801_c3_b0c0_uxn_opcodes_h_l1801_c3_b0c0_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- n8_MUX[uxn_opcodes_h_l1808_c7_e477] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1808_c7_e477_cond <= VAR_n8_MUX_uxn_opcodes_h_l1808_c7_e477_cond;
     n8_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue;
     n8_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1808_c7_e477_return_output := n8_MUX_uxn_opcodes_h_l1808_c7_e477_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1811_c7_760f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_return_output;

     -- t8_MUX[uxn_opcodes_h_l1805_c7_517b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1805_c7_517b_cond <= VAR_t8_MUX_uxn_opcodes_h_l1805_c7_517b_cond;
     t8_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue;
     t8_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1805_c7_517b_return_output := t8_MUX_uxn_opcodes_h_l1805_c7_517b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1811_c7_760f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1808_c7_e477] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1808_c7_e477_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_760f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_760f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_760f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_e477_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_e477_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_760f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1805_c7_517b_return_output;
     -- t8_MUX[uxn_opcodes_h_l1800_c2_414f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1800_c2_414f_cond <= VAR_t8_MUX_uxn_opcodes_h_l1800_c2_414f_cond;
     t8_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue;
     t8_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1800_c2_414f_return_output := t8_MUX_uxn_opcodes_h_l1800_c2_414f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1808_c7_e477] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1808_c7_e477] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1805_c7_517b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1808_c7_e477] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1805_c7_517b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1808_c7_e477] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_return_output := result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_return_output;

     -- n8_MUX[uxn_opcodes_h_l1805_c7_517b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1805_c7_517b_cond <= VAR_n8_MUX_uxn_opcodes_h_l1805_c7_517b_cond;
     n8_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue;
     n8_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1805_c7_517b_return_output := n8_MUX_uxn_opcodes_h_l1805_c7_517b_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1805_c7_517b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_e477_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_e477_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_e477_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_517b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_517b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_e477_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1800_c2_414f_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1805_c7_517b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_return_output;

     -- n8_MUX[uxn_opcodes_h_l1800_c2_414f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1800_c2_414f_cond <= VAR_n8_MUX_uxn_opcodes_h_l1800_c2_414f_cond;
     n8_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue;
     n8_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1800_c2_414f_return_output := n8_MUX_uxn_opcodes_h_l1800_c2_414f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1800_c2_414f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1805_c7_517b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1805_c7_517b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1805_c7_517b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1800_c2_414f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1800_c2_414f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_517b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_517b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_517b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_517b_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1800_c2_414f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1800_c2_414f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1800_c2_414f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1800_c2_414f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l1796_l1825_DUPLICATE_b86c LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l1796_l1825_DUPLICATE_b86c_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_4e73(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_414f_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_414f_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_414f_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_414f_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_414f_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_414f_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l1796_l1825_DUPLICATE_b86c_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l1796_l1825_DUPLICATE_b86c_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
