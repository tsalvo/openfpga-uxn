-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 37
entity dup_0CLK_6be78140 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dup_0CLK_6be78140;
architecture arch of dup_0CLK_6be78140 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2627_c6_e95f]
signal BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2627_c1_cb20]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2627_c2_0d68]
signal t8_MUX_uxn_opcodes_h_l2627_c2_0d68_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2627_c2_0d68]
signal result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2627_c2_0d68]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2627_c2_0d68]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2627_c2_0d68]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2627_c2_0d68]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2627_c2_0d68]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output : signed(3 downto 0);

-- printf_uxn_opcodes_h_l2628_c3_5617[uxn_opcodes_h_l2628_c3_5617]
signal printf_uxn_opcodes_h_l2628_c3_5617_uxn_opcodes_h_l2628_c3_5617_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2632_c11_a2a3]
signal BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2632_c7_e385]
signal t8_MUX_uxn_opcodes_h_l2632_c7_e385_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2632_c7_e385_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2632_c7_e385]
signal result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2632_c7_e385]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2632_c7_e385]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2632_c7_e385]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2632_c7_e385]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2632_c7_e385]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2635_c11_d447]
signal BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2635_c7_6374]
signal t8_MUX_uxn_opcodes_h_l2635_c7_6374_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2635_c7_6374_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2635_c7_6374]
signal result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2635_c7_6374]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2635_c7_6374]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2635_c7_6374]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2635_c7_6374]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2635_c7_6374]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_return_output : signed(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2638_c30_2d3b]
signal sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2643_c11_2509]
signal BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2643_c7_eb6d]
signal result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2643_c7_eb6d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2643_c7_eb6d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2643_c7_eb6d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2643_c7_eb6d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2648_c11_91d2]
signal BIN_OP_EQ_uxn_opcodes_h_l2648_c11_91d2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2648_c11_91d2_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2648_c11_91d2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2648_c7_cd43]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2648_c7_cd43]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f
BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_left,
BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_right,
BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_return_output);

-- t8_MUX_uxn_opcodes_h_l2627_c2_0d68
t8_MUX_uxn_opcodes_h_l2627_c2_0d68 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2627_c2_0d68_cond,
t8_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue,
t8_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse,
t8_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68
result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_cond,
result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68
result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68
result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68
result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68
result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output);

-- printf_uxn_opcodes_h_l2628_c3_5617_uxn_opcodes_h_l2628_c3_5617
printf_uxn_opcodes_h_l2628_c3_5617_uxn_opcodes_h_l2628_c3_5617 : entity work.printf_uxn_opcodes_h_l2628_c3_5617_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2628_c3_5617_uxn_opcodes_h_l2628_c3_5617_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3
BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_left,
BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_right,
BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_return_output);

-- t8_MUX_uxn_opcodes_h_l2632_c7_e385
t8_MUX_uxn_opcodes_h_l2632_c7_e385 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2632_c7_e385_cond,
t8_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue,
t8_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse,
t8_MUX_uxn_opcodes_h_l2632_c7_e385_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385
result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_cond,
result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385
result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385
result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385
result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385
result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447
BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_left,
BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_right,
BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_return_output);

-- t8_MUX_uxn_opcodes_h_l2635_c7_6374
t8_MUX_uxn_opcodes_h_l2635_c7_6374 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2635_c7_6374_cond,
t8_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue,
t8_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse,
t8_MUX_uxn_opcodes_h_l2635_c7_6374_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374
result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_cond,
result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374
result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374
result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374
result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374
result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b
sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_ins,
sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_x,
sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_y,
sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509
BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509_left,
BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509_right,
BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d
result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond,
result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d
result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d
result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d
result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2648_c11_91d2
BIN_OP_EQ_uxn_opcodes_h_l2648_c11_91d2 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2648_c11_91d2_left,
BIN_OP_EQ_uxn_opcodes_h_l2648_c11_91d2_right,
BIN_OP_EQ_uxn_opcodes_h_l2648_c11_91d2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43
result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43
result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_return_output,
 t8_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_return_output,
 t8_MUX_uxn_opcodes_h_l2632_c7_e385_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_return_output,
 t8_MUX_uxn_opcodes_h_l2635_c7_6374_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_return_output,
 sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2648_c11_91d2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2632_c7_e385_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2627_c2_0d68_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2629_c3_9c4c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2628_c3_5617_uxn_opcodes_h_l2628_c3_5617_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2635_c7_6374_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2632_c7_e385_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2633_c3_ab61 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2635_c7_6374_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2640_c3_a7c4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2645_c3_a0a9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2643_c7_eb6d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2648_c11_91d2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2648_c11_91d2_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2648_c11_91d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2632_l2627_l2643_DUPLICATE_fdcd_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2632_l2627_l2643_DUPLICATE_7292_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2632_l2648_l2627_l2643_DUPLICATE_c485_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2632_l2635_l2627_DUPLICATE_6c58_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2632_l2648_l2635_l2643_DUPLICATE_9841_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l2623_l2653_DUPLICATE_f5cb_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2640_c3_a7c4 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2640_c3_a7c4;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2629_c3_9c4c := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2629_c3_9c4c;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2633_c3_ab61 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2633_c3_ab61;
     VAR_sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2645_c3_a0a9 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2645_c3_a0a9;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2648_c11_91d2_right := to_unsigned(4, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_iffalse := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2648_c11_91d2_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse := t8;
     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2632_l2627_l2643_DUPLICATE_fdcd LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2632_l2627_l2643_DUPLICATE_fdcd_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2632_l2648_l2627_l2643_DUPLICATE_c485 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2632_l2648_l2627_l2643_DUPLICATE_c485_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2627_c6_e95f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2635_c11_d447] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_left;
     BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_return_output := BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2648_c11_91d2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2648_c11_91d2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2648_c11_91d2_left;
     BIN_OP_EQ_uxn_opcodes_h_l2648_c11_91d2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2648_c11_91d2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2648_c11_91d2_return_output := BIN_OP_EQ_uxn_opcodes_h_l2648_c11_91d2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2632_c11_a2a3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_left;
     BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_return_output := BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2632_l2648_l2635_l2643_DUPLICATE_9841 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2632_l2648_l2635_l2643_DUPLICATE_9841_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2632_l2627_l2643_DUPLICATE_7292 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2632_l2627_l2643_DUPLICATE_7292_return_output := result.is_sp_shift;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2643_c7_eb6d] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2643_c7_eb6d_return_output := result.stack_address_sp_offset;

     -- sp_relative_shift[uxn_opcodes_h_l2638_c30_2d3b] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_ins;
     sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_x;
     sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_return_output := sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2643_c11_2509] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509_left;
     BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509_return_output := BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2632_l2635_l2627_DUPLICATE_6c58 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2632_l2635_l2627_DUPLICATE_6c58_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2627_c2_0d68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2627_c6_e95f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2632_c7_e385_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_a2a3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2635_c7_6374_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2635_c11_d447_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_2509_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2648_c11_91d2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2648_c11_91d2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2632_l2635_l2627_DUPLICATE_6c58_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2632_l2635_l2627_DUPLICATE_6c58_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2632_l2635_l2627_DUPLICATE_6c58_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2632_l2648_l2635_l2643_DUPLICATE_9841_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2632_l2648_l2635_l2643_DUPLICATE_9841_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2632_l2648_l2635_l2643_DUPLICATE_9841_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2632_l2648_l2635_l2643_DUPLICATE_9841_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2632_l2627_l2643_DUPLICATE_7292_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2632_l2627_l2643_DUPLICATE_7292_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2632_l2627_l2643_DUPLICATE_7292_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2632_l2648_l2627_l2643_DUPLICATE_c485_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2632_l2648_l2627_l2643_DUPLICATE_c485_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2632_l2648_l2627_l2643_DUPLICATE_c485_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2632_l2648_l2627_l2643_DUPLICATE_c485_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2632_l2627_l2643_DUPLICATE_fdcd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2632_l2627_l2643_DUPLICATE_fdcd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2632_l2627_l2643_DUPLICATE_fdcd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2643_c7_eb6d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2638_c30_2d3b_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2648_c7_cd43] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2643_c7_eb6d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2627_c1_cb20] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2643_c7_eb6d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output := result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output;

     -- t8_MUX[uxn_opcodes_h_l2635_c7_6374] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2635_c7_6374_cond <= VAR_t8_MUX_uxn_opcodes_h_l2635_c7_6374_cond;
     t8_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue;
     t8_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2635_c7_6374_return_output := t8_MUX_uxn_opcodes_h_l2635_c7_6374_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2643_c7_eb6d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2635_c7_6374] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2648_c7_cd43] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l2628_c3_5617_uxn_opcodes_h_l2628_c3_5617_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2627_c1_cb20_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2648_c7_cd43_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2648_c7_cd43_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2635_c7_6374_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2635_c7_6374_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2635_c7_6374] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2635_c7_6374] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_return_output := result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2643_c7_eb6d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2635_c7_6374] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2643_c7_eb6d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2632_c7_e385] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_return_output;

     -- printf_uxn_opcodes_h_l2628_c3_5617[uxn_opcodes_h_l2628_c3_5617] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2628_c3_5617_uxn_opcodes_h_l2628_c3_5617_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2628_c3_5617_uxn_opcodes_h_l2628_c3_5617_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- t8_MUX[uxn_opcodes_h_l2632_c7_e385] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2632_c7_e385_cond <= VAR_t8_MUX_uxn_opcodes_h_l2632_c7_e385_cond;
     t8_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue;
     t8_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2632_c7_e385_return_output := t8_MUX_uxn_opcodes_h_l2632_c7_e385_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2635_c7_6374_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2643_c7_eb6d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2632_c7_e385_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2635_c7_6374_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2635_c7_6374_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2632_c7_e385_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2635_c7_6374] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2627_c2_0d68] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2632_c7_e385] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2632_c7_e385] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_return_output := result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_return_output;

     -- t8_MUX[uxn_opcodes_h_l2627_c2_0d68] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2627_c2_0d68_cond <= VAR_t8_MUX_uxn_opcodes_h_l2627_c2_0d68_cond;
     t8_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue;
     t8_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output := t8_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2635_c7_6374] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2632_c7_e385] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2635_c7_6374_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_e385_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2635_c7_6374_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_e385_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_e385_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2627_c2_0d68] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2632_c7_e385] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2627_c2_0d68] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2632_c7_e385] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2627_c2_0d68] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output := result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_e385_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_e385_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2627_c2_0d68] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2627_c2_0d68] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l2623_l2653_DUPLICATE_f5cb LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l2623_l2653_DUPLICATE_f5cb_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2627_c2_0d68_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l2623_l2653_DUPLICATE_f5cb_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l2623_l2653_DUPLICATE_f5cb_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
