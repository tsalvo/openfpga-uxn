-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 36
entity nip2_0CLK_1a2ef46d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end nip2_0CLK_1a2ef46d;
architecture arch of nip2_0CLK_1a2ef46d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2174_c6_2905]
signal BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2174_c2_d609]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2174_c2_d609]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2174_c2_d609]
signal result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2174_c2_d609]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2174_c2_d609]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2174_c2_d609]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2174_c2_d609]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_return_output : unsigned(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2174_c2_d609]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2174_c2_d609]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2174_c2_d609]
signal t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2174_c2_d609]
signal t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2187_c11_d5c4]
signal BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2187_c7_40d4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2187_c7_40d4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2187_c7_40d4]
signal result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2187_c7_40d4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2187_c7_40d4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2187_c7_40d4]
signal t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2187_c7_40d4]
signal t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2190_c11_d11e]
signal BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2190_c7_6598]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2190_c7_6598]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2190_c7_6598]
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2190_c7_6598]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2190_c7_6598]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2190_c7_6598]
signal t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2190_c7_6598]
signal t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2192_c30_b2a0]
signal sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2197_c11_3ef4]
signal BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2197_c7_1d10]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2197_c7_1d10]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2197_c7_1d10]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2197_c7_1d10]
signal result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output : unsigned(7 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2197_c7_1d10]
signal t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_pc_updated := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.is_ram_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;
      base.is_stack_index_flipped := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905
BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_left,
BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_right,
BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609
result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609
result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609
result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_cond,
result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609
result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609
result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609
result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609
result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2174_c2_d609
t16_low_MUX_uxn_opcodes_h_l2174_c2_d609 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_cond,
t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue,
t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse,
t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2174_c2_d609
t16_high_MUX_uxn_opcodes_h_l2174_c2_d609 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_cond,
t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue,
t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse,
t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4
BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_left,
BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_right,
BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_cond,
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4
t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_cond,
t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue,
t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse,
t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4
t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_cond,
t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue,
t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse,
t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e
BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_left,
BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_right,
BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_cond,
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2190_c7_6598
t16_low_MUX_uxn_opcodes_h_l2190_c7_6598 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_cond,
t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue,
t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse,
t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2190_c7_6598
t16_high_MUX_uxn_opcodes_h_l2190_c7_6598 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_cond,
t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue,
t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse,
t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0
sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_ins,
sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_x,
sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_y,
sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4
BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4_left,
BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4_right,
BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_cond,
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10
t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_cond,
t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue,
t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse,
t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_return_output,
 t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_return_output,
 t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output,
 t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output,
 t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_return_output,
 t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_return_output,
 t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_return_output,
 sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output,
 t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2174_c2_d609_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2174_c2_d609_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2174_c2_d609_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2179_c3_5c52 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2184_c3_ffa4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2174_c2_d609_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2188_c3_85a3 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2194_c3_8d3b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2200_c3_7ab6 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2197_c7_1d10_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2199_c3_f37c : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2174_l2197_l2187_DUPLICATE_c410_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2197_l2187_DUPLICATE_d39f_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_9121_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2197_l2187_l2190_DUPLICATE_a49d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l2205_l2170_DUPLICATE_7344_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2200_c3_7ab6 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2200_c3_7ab6;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2194_c3_8d3b := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2194_c3_8d3b;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2199_c3_f37c := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2199_c3_f37c;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2188_c3_85a3 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2188_c3_85a3;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2184_c3_ffa4 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2184_c3_ffa4;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2179_c3_5c52 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2179_c3_5c52;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_y := resize(to_signed(-2, 3), 4);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue := VAR_previous_stack_read;
     VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse := t16_high;
     VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse := t16_low;
     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2174_c2_d609] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2174_c2_d609_return_output := result.is_vram_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2197_l2187_DUPLICATE_d39f LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2197_l2187_DUPLICATE_d39f_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2197_l2187_l2190_DUPLICATE_a49d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2197_l2187_l2190_DUPLICATE_a49d_return_output := result.is_opc_done;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2174_c2_d609] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2174_c2_d609_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l2174_c6_2905] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_left;
     BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_return_output := BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2192_c30_b2a0] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_ins;
     sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_x;
     sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_return_output := sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2174_c2_d609] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2174_c2_d609_return_output := result.is_ram_write;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2197_c7_1d10] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2197_c7_1d10_return_output := result.stack_address_sp_offset;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2174_c2_d609] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2174_c2_d609_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_9121 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_9121_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2187_c11_d5c4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_left;
     BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_return_output := BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2197_c11_3ef4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4_left;
     BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4_return_output := BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2174_l2197_l2187_DUPLICATE_c410 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2174_l2197_l2187_DUPLICATE_c410_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2190_c11_d11e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_2905_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_d5c4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_d11e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_3ef4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2197_l2187_DUPLICATE_d39f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2197_l2187_DUPLICATE_d39f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2197_l2187_l2190_DUPLICATE_a49d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2197_l2187_l2190_DUPLICATE_a49d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2197_l2187_l2190_DUPLICATE_a49d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_9121_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_9121_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2174_l2197_l2187_DUPLICATE_c410_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2174_l2197_l2187_DUPLICATE_c410_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2174_l2197_l2187_DUPLICATE_c410_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2174_c2_d609_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2174_c2_d609_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2174_c2_d609_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2174_c2_d609_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2197_c7_1d10_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_b2a0_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2197_c7_1d10] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output := result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2190_c7_6598] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2174_c2_d609] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2197_c7_1d10] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2174_c2_d609] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2174_c2_d609] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2190_c7_6598] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_cond;
     t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_return_output := t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2197_c7_1d10] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2174_c2_d609] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2197_c7_1d10] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2197_c7_1d10] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_cond;
     t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output := t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_6598_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_6598_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_1d10_return_output;
     -- t16_high_MUX[uxn_opcodes_h_l2187_c7_40d4] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_cond;
     t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output := t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2190_c7_6598] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2190_c7_6598] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2187_c7_40d4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2190_c7_6598] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_cond;
     t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_return_output := t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2190_c7_6598] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_return_output := result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2190_c7_6598] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_6598_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_6598_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_6598_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_6598_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_6598_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2187_c7_40d4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2174_c2_d609] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_cond;
     t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_return_output := t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2187_c7_40d4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2174_c2_d609] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2187_c7_40d4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output := result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2187_c7_40d4] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_cond;
     t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output := t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2187_c7_40d4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output;
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_d609_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_40d4_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2174_c2_d609] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2174_c2_d609] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_cond;
     t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_return_output := t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2174_c2_d609] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2174_c2_d609] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_return_output := result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2174_c2_d609] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_return_output;

     -- Submodule level 5
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_d609_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l2205_l2170_DUPLICATE_7344 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l2205_l2170_DUPLICATE_7344_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6(
     result,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_d609_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_d609_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_d609_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_d609_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_d609_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_d609_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_d609_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_d609_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_d609_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l2205_l2170_DUPLICATE_7344_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l2205_l2170_DUPLICATE_7344_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
