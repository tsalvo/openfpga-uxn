-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 52
entity ldr_0CLK_c61094da is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldr_0CLK_c61094da;
architecture arch of ldr_0CLK_c61094da is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1524_c6_18e1]
signal BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1524_c1_08e3]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1524_c2_5b97]
signal t8_MUX_uxn_opcodes_h_l1524_c2_5b97_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1524_c2_5b97]
signal result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1524_c2_5b97]
signal result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1524_c2_5b97]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1524_c2_5b97]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1524_c2_5b97]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1524_c2_5b97]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1524_c2_5b97]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output : signed(3 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1524_c2_5b97]
signal tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1525_c3_9e70[uxn_opcodes_h_l1525_c3_9e70]
signal printf_uxn_opcodes_h_l1525_c3_9e70_uxn_opcodes_h_l1525_c3_9e70_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1529_c11_a626]
signal BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1529_c7_17e5]
signal t8_MUX_uxn_opcodes_h_l1529_c7_17e5_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1529_c7_17e5]
signal result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1529_c7_17e5]
signal result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1529_c7_17e5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1529_c7_17e5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1529_c7_17e5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1529_c7_17e5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1529_c7_17e5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output : signed(3 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1529_c7_17e5]
signal tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1532_c11_24ec]
signal BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1532_c7_65bc]
signal t8_MUX_uxn_opcodes_h_l1532_c7_65bc_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1532_c7_65bc]
signal result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1532_c7_65bc]
signal result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1532_c7_65bc]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1532_c7_65bc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1532_c7_65bc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1532_c7_65bc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1532_c7_65bc]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output : signed(3 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1532_c7_65bc]
signal tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1535_c30_a1c1]
signal sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_return_output : signed(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1536_c22_7deb]
signal BIN_OP_PLUS_uxn_opcodes_h_l1536_c22_7deb_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1536_c22_7deb_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1536_c22_7deb_return_output : signed(17 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1538_c11_d9e0]
signal BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1538_c7_36a4]
signal result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1538_c7_36a4]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1538_c7_36a4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1538_c7_36a4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1538_c7_36a4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output : unsigned(3 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1538_c7_36a4]
signal tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1541_c11_81c2]
signal BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1541_c7_1446]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1541_c7_1446]
signal result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1541_c7_1446]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1541_c7_1446]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1541_c7_1446]
signal tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1547_c11_5e96]
signal BIN_OP_EQ_uxn_opcodes_h_l1547_c11_5e96_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1547_c11_5e96_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1547_c11_5e96_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1547_c7_b9a0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1547_c7_b9a0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_return_output : unsigned(0 downto 0);

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_a310( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u16_value := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1
BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_left,
BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_right,
BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_return_output);

-- t8_MUX_uxn_opcodes_h_l1524_c2_5b97
t8_MUX_uxn_opcodes_h_l1524_c2_5b97 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1524_c2_5b97_cond,
t8_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue,
t8_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse,
t8_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97
result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_cond,
result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97
result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_cond,
result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97
result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97
result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97
result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97
result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97
tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_cond,
tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue,
tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse,
tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output);

-- printf_uxn_opcodes_h_l1525_c3_9e70_uxn_opcodes_h_l1525_c3_9e70
printf_uxn_opcodes_h_l1525_c3_9e70_uxn_opcodes_h_l1525_c3_9e70 : entity work.printf_uxn_opcodes_h_l1525_c3_9e70_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1525_c3_9e70_uxn_opcodes_h_l1525_c3_9e70_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626
BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_left,
BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_right,
BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_return_output);

-- t8_MUX_uxn_opcodes_h_l1529_c7_17e5
t8_MUX_uxn_opcodes_h_l1529_c7_17e5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1529_c7_17e5_cond,
t8_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue,
t8_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse,
t8_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5
result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_cond,
result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5
result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_cond,
result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5
result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5
result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5
result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5
result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5
tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_cond,
tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue,
tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse,
tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec
BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_left,
BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_right,
BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_return_output);

-- t8_MUX_uxn_opcodes_h_l1532_c7_65bc
t8_MUX_uxn_opcodes_h_l1532_c7_65bc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1532_c7_65bc_cond,
t8_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue,
t8_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse,
t8_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc
result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_cond,
result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc
result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_cond,
result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc
result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc
result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc
result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc
result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc
tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_cond,
tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue,
tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse,
tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1
sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_ins,
sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_x,
sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_y,
sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1536_c22_7deb
BIN_OP_PLUS_uxn_opcodes_h_l1536_c22_7deb : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1536_c22_7deb_left,
BIN_OP_PLUS_uxn_opcodes_h_l1536_c22_7deb_right,
BIN_OP_PLUS_uxn_opcodes_h_l1536_c22_7deb_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0
BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0_left,
BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0_right,
BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4
result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_cond,
result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4
result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4
result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4
result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4
tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_cond,
tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue,
tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse,
tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2
BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2_left,
BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2_right,
BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446
result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_cond,
result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446
result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446
result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1541_c7_1446
tmp8_MUX_uxn_opcodes_h_l1541_c7_1446 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_cond,
tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue,
tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse,
tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1547_c11_5e96
BIN_OP_EQ_uxn_opcodes_h_l1547_c11_5e96 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1547_c11_5e96_left,
BIN_OP_EQ_uxn_opcodes_h_l1547_c11_5e96_right,
BIN_OP_EQ_uxn_opcodes_h_l1547_c11_5e96_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0
result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0
result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_return_output,
 t8_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output,
 tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_return_output,
 t8_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output,
 tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_return_output,
 t8_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output,
 tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output,
 sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1536_c22_7deb_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output,
 tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_return_output,
 tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1547_c11_5e96_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1524_c2_5b97_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1526_c3_8f2f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1525_c3_9e70_uxn_opcodes_h_l1525_c3_9e70_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1529_c7_17e5_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1530_c3_4703 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1532_c7_65bc_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l1536_c3_c133 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1536_c22_7deb_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l1536_c27_336c_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1536_c22_7deb_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1536_c22_7deb_return_output : signed(17 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1544_c3_d340 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1547_c11_5e96_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1547_c11_5e96_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1547_c11_5e96_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1529_l1532_l1524_DUPLICATE_a968_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1541_l1538_l1532_l1529_l1524_DUPLICATE_2285_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1529_l1524_l1538_DUPLICATE_c100_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1538_l1532_l1529_l1524_l1547_DUPLICATE_e1be_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1529_l1532_l1524_DUPLICATE_c052_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1541_l1538_l1532_l1529_l1547_DUPLICATE_55d4_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1541_l1532_l1538_DUPLICATE_8568_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a310_uxn_opcodes_h_l1520_l1552_DUPLICATE_e614_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1530_c3_4703 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1530_c3_4703;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1526_c3_8f2f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1526_c3_8f2f;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1544_c3_d340 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1544_c3_d340;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1547_c11_5e96_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_right := to_unsigned(2, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_ins := VAR_ins;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1536_c22_7deb_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1547_c11_5e96_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse := tmp8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1529_l1524_l1538_DUPLICATE_c100 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1529_l1524_l1538_DUPLICATE_c100_return_output := result.is_sp_shift;

     -- sp_relative_shift[uxn_opcodes_h_l1535_c30_a1c1] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_ins;
     sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_x;
     sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_return_output := sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1532_c11_24ec] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_left;
     BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_return_output := BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_return_output;

     -- CAST_TO_int8_t[uxn_opcodes_h_l1536_c27_336c] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l1536_c27_336c_return_output := CAST_TO_int8_t_uint8_t(
     VAR_previous_stack_read);

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1529_l1532_l1524_DUPLICATE_c052 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1529_l1532_l1524_DUPLICATE_c052_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1529_l1532_l1524_DUPLICATE_a968 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1529_l1532_l1524_DUPLICATE_a968_return_output := result.u16_value;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1541_l1532_l1538_DUPLICATE_8568 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1541_l1532_l1538_DUPLICATE_8568_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1524_c6_18e1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_left;
     BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_return_output := BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1541_l1538_l1532_l1529_l1524_DUPLICATE_2285 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1541_l1538_l1532_l1529_l1524_DUPLICATE_2285_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1541_l1538_l1532_l1529_l1547_DUPLICATE_55d4 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1541_l1538_l1532_l1529_l1547_DUPLICATE_55d4_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1538_l1532_l1529_l1524_l1547_DUPLICATE_e1be LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1538_l1532_l1529_l1524_l1547_DUPLICATE_e1be_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1541_c11_81c2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2_left;
     BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2_return_output := BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1547_c11_5e96] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1547_c11_5e96_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1547_c11_5e96_left;
     BIN_OP_EQ_uxn_opcodes_h_l1547_c11_5e96_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1547_c11_5e96_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1547_c11_5e96_return_output := BIN_OP_EQ_uxn_opcodes_h_l1547_c11_5e96_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1538_c11_d9e0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0_left;
     BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0_return_output := BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1529_c11_a626] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_left;
     BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_return_output := BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1524_c2_5b97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1524_c6_18e1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1529_c7_17e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1529_c11_a626_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1532_c7_65bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_24ec_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1538_c11_d9e0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1541_c11_81c2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1547_c11_5e96_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1547_c11_5e96_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1536_c22_7deb_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l1536_c27_336c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1529_l1532_l1524_DUPLICATE_c052_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1529_l1532_l1524_DUPLICATE_c052_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1529_l1532_l1524_DUPLICATE_c052_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1529_l1532_l1524_DUPLICATE_a968_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1529_l1532_l1524_DUPLICATE_a968_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1529_l1532_l1524_DUPLICATE_a968_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1541_l1538_l1532_l1529_l1547_DUPLICATE_55d4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1541_l1538_l1532_l1529_l1547_DUPLICATE_55d4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1541_l1538_l1532_l1529_l1547_DUPLICATE_55d4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1541_l1538_l1532_l1529_l1547_DUPLICATE_55d4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1541_l1538_l1532_l1529_l1547_DUPLICATE_55d4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1529_l1524_l1538_DUPLICATE_c100_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1529_l1524_l1538_DUPLICATE_c100_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1529_l1524_l1538_DUPLICATE_c100_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1538_l1532_l1529_l1524_l1547_DUPLICATE_e1be_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1538_l1532_l1529_l1524_l1547_DUPLICATE_e1be_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1538_l1532_l1529_l1524_l1547_DUPLICATE_e1be_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1538_l1532_l1529_l1524_l1547_DUPLICATE_e1be_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1538_l1532_l1529_l1524_l1547_DUPLICATE_e1be_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1541_l1532_l1538_DUPLICATE_8568_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1541_l1532_l1538_DUPLICATE_8568_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1541_l1532_l1538_DUPLICATE_8568_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1541_l1538_l1532_l1529_l1524_DUPLICATE_2285_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1541_l1538_l1532_l1529_l1524_DUPLICATE_2285_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1541_l1538_l1532_l1529_l1524_DUPLICATE_2285_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1541_l1538_l1532_l1529_l1524_DUPLICATE_2285_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1541_l1538_l1532_l1529_l1524_DUPLICATE_2285_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1535_c30_a1c1_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1541_c7_1446] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_return_output := result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_return_output;

     -- t8_MUX[uxn_opcodes_h_l1532_c7_65bc] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1532_c7_65bc_cond <= VAR_t8_MUX_uxn_opcodes_h_l1532_c7_65bc_cond;
     t8_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue;
     t8_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output := t8_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1532_c7_65bc] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1547_c7_b9a0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1538_c7_36a4] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1541_c7_1446] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_cond;
     tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_return_output := tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1536_c22_7deb] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1536_c22_7deb_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1536_c22_7deb_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1536_c22_7deb_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1536_c22_7deb_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1536_c22_7deb_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1536_c22_7deb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1541_c7_1446] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1547_c7_b9a0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1524_c1_08e3] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_return_output;

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l1536_c3_c133 := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1536_c22_7deb_return_output)),16);
     VAR_printf_uxn_opcodes_h_l1525_c3_9e70_uxn_opcodes_h_l1525_c3_9e70_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1524_c1_08e3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1547_c7_b9a0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1547_c7_b9a0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1541_c7_1446_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1541_c7_1446_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1541_c7_1446_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue := VAR_result_u16_value_uxn_opcodes_h_l1536_c3_c133;
     -- t8_MUX[uxn_opcodes_h_l1529_c7_17e5] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1529_c7_17e5_cond <= VAR_t8_MUX_uxn_opcodes_h_l1529_c7_17e5_cond;
     t8_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue;
     t8_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output := t8_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1529_c7_17e5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1532_c7_65bc] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output := result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1538_c7_36a4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output := result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1532_c7_65bc] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1538_c7_36a4] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_cond;
     tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output := tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1541_c7_1446] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_return_output;

     -- printf_uxn_opcodes_h_l1525_c3_9e70[uxn_opcodes_h_l1525_c3_9e70] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1525_c3_9e70_uxn_opcodes_h_l1525_c3_9e70_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1525_c3_9e70_uxn_opcodes_h_l1525_c3_9e70_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1538_c7_36a4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1541_c7_1446] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1541_c7_1446_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1541_c7_1446_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1529_c7_17e5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output;

     -- t8_MUX[uxn_opcodes_h_l1524_c2_5b97] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1524_c2_5b97_cond <= VAR_t8_MUX_uxn_opcodes_h_l1524_c2_5b97_cond;
     t8_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue;
     t8_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output := t8_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1538_c7_36a4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1529_c7_17e5] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output := result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1532_c7_65bc] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output := result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1524_c2_5b97] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1532_c7_65bc] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_cond;
     tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output := tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1538_c7_36a4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1532_c7_65bc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1538_c7_36a4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l1524_c2_5b97] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output := result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1524_c2_5b97] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1529_c7_17e5] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_cond;
     tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output := tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1529_c7_17e5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1529_c7_17e5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output := result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1532_c7_65bc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1532_c7_65bc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_65bc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1529_c7_17e5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1529_c7_17e5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1524_c2_5b97] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_cond;
     tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output := tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1524_c2_5b97] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output := result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1524_c2_5b97] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1529_c7_17e5_return_output;
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1524_c2_5b97] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1524_c2_5b97] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a310_uxn_opcodes_h_l1520_l1552_DUPLICATE_e614 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a310_uxn_opcodes_h_l1520_l1552_DUPLICATE_e614_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a310(
     result,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1524_c2_5b97_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a310_uxn_opcodes_h_l1520_l1552_DUPLICATE_e614_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a310_uxn_opcodes_h_l1520_l1552_DUPLICATE_e614_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
