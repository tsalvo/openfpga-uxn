-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 47
entity ldz_0CLK_b128164d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldz_0CLK_b128164d;
architecture arch of ldz_0CLK_b128164d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1454_c6_6169]
signal BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1454_c2_0e60]
signal tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1454_c2_0e60]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1454_c2_0e60]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1454_c2_0e60]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1454_c2_0e60]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1454_c2_0e60]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1454_c2_0e60]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1454_c2_0e60]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1454_c2_0e60]
signal result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1454_c2_0e60]
signal result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(7 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1454_c2_0e60]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1454_c2_0e60]
signal t8_MUX_uxn_opcodes_h_l1454_c2_0e60_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1467_c11_b2a3]
signal BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1467_c7_4c24]
signal tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1467_c7_4c24]
signal result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1467_c7_4c24]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1467_c7_4c24]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1467_c7_4c24]
signal result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1467_c7_4c24]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1467_c7_4c24]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1467_c7_4c24]
signal t8_MUX_uxn_opcodes_h_l1467_c7_4c24_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1470_c11_00f8]
signal BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1470_c7_7f6c]
signal tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1470_c7_7f6c]
signal result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1470_c7_7f6c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1470_c7_7f6c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1470_c7_7f6c]
signal result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1470_c7_7f6c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1470_c7_7f6c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1470_c7_7f6c]
signal t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1472_c30_c692]
signal sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1475_c11_9abb]
signal BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1475_c7_c176]
signal tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1475_c7_c176]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1475_c7_c176]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1475_c7_c176]
signal result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1475_c7_c176]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1475_c7_c176]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1478_c11_2878]
signal BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1478_c7_4acb]
signal tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1478_c7_4acb]
signal result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1478_c7_4acb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1478_c7_4acb]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1478_c7_4acb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output : unsigned(3 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_42c1( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_ram_write := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_index_flipped := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.u16_value := ref_toks_8;
      base.u8_value := ref_toks_9;
      base.is_vram_write := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169
BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_left,
BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_right,
BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60
tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_cond,
tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue,
tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse,
tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60
result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60
result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60
result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60
result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60
result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60
result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_cond,
result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60
result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_cond,
result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60
result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output);

-- t8_MUX_uxn_opcodes_h_l1454_c2_0e60
t8_MUX_uxn_opcodes_h_l1454_c2_0e60 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1454_c2_0e60_cond,
t8_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue,
t8_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse,
t8_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3
BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_left,
BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_right,
BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24
tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_cond,
tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue,
tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse,
tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24
result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_cond,
result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24
result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24
result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24
result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_cond,
result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24
result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output);

-- t8_MUX_uxn_opcodes_h_l1467_c7_4c24
t8_MUX_uxn_opcodes_h_l1467_c7_4c24 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1467_c7_4c24_cond,
t8_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue,
t8_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse,
t8_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8
BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_left,
BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_right,
BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c
tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond,
tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue,
tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse,
tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c
result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond,
result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c
result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c
result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c
result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c
result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output);

-- t8_MUX_uxn_opcodes_h_l1470_c7_7f6c
t8_MUX_uxn_opcodes_h_l1470_c7_7f6c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond,
t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue,
t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse,
t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1472_c30_c692
sp_relative_shift_uxn_opcodes_h_l1472_c30_c692 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_ins,
sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_x,
sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_y,
sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb
BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb_left,
BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb_right,
BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1475_c7_c176
tmp8_MUX_uxn_opcodes_h_l1475_c7_c176 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_cond,
tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue,
tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse,
tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176
result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176
result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176
result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_cond,
result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176
result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878
BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878_left,
BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878_right,
BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb
tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_cond,
tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue,
tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse,
tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb
result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_cond,
result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb
result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb
result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_return_output,
 tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output,
 t8_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_return_output,
 tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output,
 t8_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_return_output,
 tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output,
 t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output,
 sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb_return_output,
 tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878_return_output,
 tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1459_c3_ddde : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1464_c3_eaba : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1454_c2_0e60_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1468_c3_6844 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1467_c7_4c24_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1473_c22_1f3e_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1476_c3_2983 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1481_c3_493f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1454_l1467_l1470_DUPLICATE_90ab_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1478_l1475_l1470_l1467_l1454_DUPLICATE_0f92_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1475_l1467_l1478_l1470_DUPLICATE_9c23_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1475_l1467_DUPLICATE_d0de_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1475_l1467_l1478_l1470_DUPLICATE_9574_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1475_l1478_l1470_DUPLICATE_6771_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_42c1_uxn_opcodes_h_l1486_l1450_DUPLICATE_a91a_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_right := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1476_c3_2983 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1476_c3_2983;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1481_c3_493f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1481_c3_493f;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1464_c3_eaba := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1464_c3_eaba;
     VAR_sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_right := to_unsigned(2, 2);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1468_c3_6844 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1468_c3_6844;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1459_c3_ddde := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1459_c3_ddde;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse := tmp8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1470_c11_00f8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_left;
     BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_return_output := BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1454_c6_6169] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_left;
     BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_return_output := BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1467_c11_b2a3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_left;
     BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_return_output := BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1472_c30_c692] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_ins;
     sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_x;
     sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_return_output := sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1454_l1467_l1470_DUPLICATE_90ab LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1454_l1467_l1470_DUPLICATE_90ab_return_output := result.u16_value;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1454_c2_0e60] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1454_c2_0e60_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1475_l1467_l1478_l1470_DUPLICATE_9c23 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1475_l1467_l1478_l1470_DUPLICATE_9c23_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1475_l1478_l1470_DUPLICATE_6771 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1475_l1478_l1470_DUPLICATE_6771_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1475_c11_9abb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb_left;
     BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb_return_output := BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1478_l1475_l1470_l1467_l1454_DUPLICATE_0f92 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1478_l1475_l1470_l1467_l1454_DUPLICATE_0f92_return_output := result.u8_value;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1454_c2_0e60] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1454_c2_0e60_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l1478_c11_2878] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878_left;
     BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878_return_output := BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1475_l1467_DUPLICATE_d0de LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1475_l1467_DUPLICATE_d0de_return_output := result.sp_relative_shift;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1454_c2_0e60] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1454_c2_0e60_return_output := result.is_vram_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1454_c2_0e60] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1454_c2_0e60_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1475_l1467_l1478_l1470_DUPLICATE_9574 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1475_l1467_l1478_l1470_DUPLICATE_9574_return_output := result.is_stack_write;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1473_c22_1f3e] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1473_c22_1f3e_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1454_c2_0e60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1454_c6_6169_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1467_c7_4c24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1467_c11_b2a3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1470_c11_00f8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1475_c11_9abb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1478_c11_2878_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1473_c22_1f3e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1475_l1467_DUPLICATE_d0de_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1475_l1467_DUPLICATE_d0de_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1454_l1467_l1470_DUPLICATE_90ab_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1454_l1467_l1470_DUPLICATE_90ab_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1454_l1467_l1470_DUPLICATE_90ab_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1475_l1467_l1478_l1470_DUPLICATE_9c23_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1475_l1467_l1478_l1470_DUPLICATE_9c23_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1475_l1467_l1478_l1470_DUPLICATE_9c23_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1475_l1467_l1478_l1470_DUPLICATE_9c23_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1475_l1467_l1478_l1470_DUPLICATE_9574_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1475_l1467_l1478_l1470_DUPLICATE_9574_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1475_l1467_l1478_l1470_DUPLICATE_9574_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1475_l1467_l1478_l1470_DUPLICATE_9574_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1475_l1478_l1470_DUPLICATE_6771_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1475_l1478_l1470_DUPLICATE_6771_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1475_l1478_l1470_DUPLICATE_6771_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1478_l1475_l1470_l1467_l1454_DUPLICATE_0f92_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1478_l1475_l1470_l1467_l1454_DUPLICATE_0f92_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1478_l1475_l1470_l1467_l1454_DUPLICATE_0f92_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1478_l1475_l1470_l1467_l1454_DUPLICATE_0f92_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1478_l1475_l1470_l1467_l1454_DUPLICATE_0f92_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1454_c2_0e60_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1454_c2_0e60_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1454_c2_0e60_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1454_c2_0e60_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1472_c30_c692_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1454_c2_0e60] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1478_c7_4acb] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1454_c2_0e60] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1478_c7_4acb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1478_c7_4acb] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_cond;
     tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output := tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1454_c2_0e60] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1478_c7_4acb] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output := result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output;

     -- t8_MUX[uxn_opcodes_h_l1470_c7_7f6c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond <= VAR_t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond;
     t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue;
     t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output := t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1454_c2_0e60] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1478_c7_4acb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1470_c7_7f6c] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output := result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1475_c7_c176] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1475_c7_c176_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1478_c7_4acb_return_output;
     -- t8_MUX[uxn_opcodes_h_l1467_c7_4c24] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1467_c7_4c24_cond <= VAR_t8_MUX_uxn_opcodes_h_l1467_c7_4c24_cond;
     t8_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue;
     t8_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output := t8_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1470_c7_7f6c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1475_c7_c176] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_cond;
     tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_return_output := tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1475_c7_c176] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1475_c7_c176] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_return_output := result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1467_c7_4c24] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output := result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1475_c7_c176] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1475_c7_c176] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1475_c7_c176_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1475_c7_c176_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1475_c7_c176_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1475_c7_c176_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1475_c7_c176_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l1454_c2_0e60] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output := result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1470_c7_7f6c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1470_c7_7f6c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1470_c7_7f6c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1470_c7_7f6c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1467_c7_4c24] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1470_c7_7f6c] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_cond;
     tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output := tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output;

     -- t8_MUX[uxn_opcodes_h_l1454_c2_0e60] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1454_c2_0e60_cond <= VAR_t8_MUX_uxn_opcodes_h_l1454_c2_0e60_cond;
     t8_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue;
     t8_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output := t8_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1470_c7_7f6c_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1467_c7_4c24] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1467_c7_4c24] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output := result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1454_c2_0e60] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1467_c7_4c24] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_cond;
     tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output := tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1467_c7_4c24] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1467_c7_4c24] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1467_c7_4c24_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1454_c2_0e60] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1454_c2_0e60] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1454_c2_0e60] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output := result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1454_c2_0e60] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_cond;
     tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output := tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1454_c2_0e60] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output;

     -- Submodule level 6
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_42c1_uxn_opcodes_h_l1486_l1450_DUPLICATE_a91a LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_42c1_uxn_opcodes_h_l1486_l1450_DUPLICATE_a91a_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_42c1(
     result,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1454_c2_0e60_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_42c1_uxn_opcodes_h_l1486_l1450_DUPLICATE_a91a_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_42c1_uxn_opcodes_h_l1486_l1450_DUPLICATE_a91a_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
