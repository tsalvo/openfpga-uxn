-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 33
entity VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_0CLK_6481cb28 is
port(
 elem_val : in unsigned(7 downto 0);
 ref_toks_0 : in uint8_t_16;
 var_dim_0 : in unsigned(3 downto 0);
 return_output : out uint8_t_array_16_t);
end VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_0CLK_6481cb28;
architecture arch of VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_0CLK_6481cb28 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d584]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d584_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d584_right : unsigned(1 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d584_return_output : unsigned(0 downto 0);

-- rv_data_2_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a]
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_cond : unsigned(0 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_iftrue : unsigned(7 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_iffalse : unsigned(7 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_492e]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_492e_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_492e_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_492e_return_output : unsigned(0 downto 0);

-- rv_data_8_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d]
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_cond : unsigned(0 downto 0);
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_iftrue : unsigned(7 downto 0);
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_iffalse : unsigned(7 downto 0);
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_3a2b]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_3a2b_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_3a2b_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_3a2b_return_output : unsigned(0 downto 0);

-- rv_data_5_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43]
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_cond : unsigned(0 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_iftrue : unsigned(7 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_iffalse : unsigned(7 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_8c77]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_8c77_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_8c77_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_8c77_return_output : unsigned(0 downto 0);

-- rv_data_11_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171]
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_cond : unsigned(0 downto 0);
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_iftrue : unsigned(7 downto 0);
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_iffalse : unsigned(7 downto 0);
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_8777]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_8777_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_8777_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_8777_return_output : unsigned(0 downto 0);

-- rv_data_14_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431]
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_cond : unsigned(0 downto 0);
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_iftrue : unsigned(7 downto 0);
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_iffalse : unsigned(7 downto 0);
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_493d]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_493d_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_493d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_493d_return_output : unsigned(0 downto 0);

-- rv_data_0_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c]
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_cond : unsigned(0 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_iftrue : unsigned(7 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_iffalse : unsigned(7 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_6132]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_6132_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_6132_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_6132_return_output : unsigned(0 downto 0);

-- rv_data_6_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506]
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_cond : unsigned(0 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_iftrue : unsigned(7 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_iffalse : unsigned(7 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_cc1e]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_cc1e_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_cc1e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_cc1e_return_output : unsigned(0 downto 0);

-- rv_data_3_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8]
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_cond : unsigned(0 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_iftrue : unsigned(7 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_iffalse : unsigned(7 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_9d6a]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_9d6a_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_9d6a_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_9d6a_return_output : unsigned(0 downto 0);

-- rv_data_9_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea]
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_cond : unsigned(0 downto 0);
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_iftrue : unsigned(7 downto 0);
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_iffalse : unsigned(7 downto 0);
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_8a43]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_8a43_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_8a43_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_8a43_return_output : unsigned(0 downto 0);

-- rv_data_15_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c]
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_cond : unsigned(0 downto 0);
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_iftrue : unsigned(7 downto 0);
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_iffalse : unsigned(7 downto 0);
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_814e]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_814e_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_814e_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_814e_return_output : unsigned(0 downto 0);

-- rv_data_12_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3]
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_cond : unsigned(0 downto 0);
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_iftrue : unsigned(7 downto 0);
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_iffalse : unsigned(7 downto 0);
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_84b5]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_84b5_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_84b5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_84b5_return_output : unsigned(0 downto 0);

-- rv_data_1_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d]
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_cond : unsigned(0 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_iftrue : unsigned(7 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_iffalse : unsigned(7 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_577e]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_577e_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_577e_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_577e_return_output : unsigned(0 downto 0);

-- rv_data_4_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741]
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_cond : unsigned(0 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_iftrue : unsigned(7 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_iffalse : unsigned(7 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_05b3]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_05b3_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_05b3_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_05b3_return_output : unsigned(0 downto 0);

-- rv_data_7_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778]
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_cond : unsigned(0 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_iftrue : unsigned(7 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_iffalse : unsigned(7 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_a903]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_a903_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_a903_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_a903_return_output : unsigned(0 downto 0);

-- rv_data_13_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b]
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_cond : unsigned(0 downto 0);
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_iftrue : unsigned(7 downto 0);
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_iffalse : unsigned(7 downto 0);
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_848c]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_848c_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_848c_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_848c_return_output : unsigned(0 downto 0);

-- rv_data_10_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf]
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_cond : unsigned(0 downto 0);
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_iftrue : unsigned(7 downto 0);
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_iffalse : unsigned(7 downto 0);
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_return_output : unsigned(7 downto 0);

function CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_eae2( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned) return uint8_t_array_16_t is
 
  variable base : uint8_t_array_16_t; 
  variable return_output : uint8_t_array_16_t;
begin
      base.data(2) := ref_toks_0;
      base.data(8) := ref_toks_1;
      base.data(5) := ref_toks_2;
      base.data(11) := ref_toks_3;
      base.data(14) := ref_toks_4;
      base.data(0) := ref_toks_5;
      base.data(6) := ref_toks_6;
      base.data(3) := ref_toks_7;
      base.data(9) := ref_toks_8;
      base.data(15) := ref_toks_9;
      base.data(12) := ref_toks_10;
      base.data(1) := ref_toks_11;
      base.data(4) := ref_toks_12;
      base.data(7) := ref_toks_13;
      base.data(13) := ref_toks_14;
      base.data(10) := ref_toks_15;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d584
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d584 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d584_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d584_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d584_return_output);

-- rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_cond,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_iftrue,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_iffalse,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_492e
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_492e : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_492e_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_492e_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_492e_return_output);

-- rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_cond,
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_iftrue,
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_iffalse,
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_3a2b
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_3a2b : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_3a2b_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_3a2b_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_3a2b_return_output);

-- rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_cond,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_iftrue,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_iffalse,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_8c77
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_8c77 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_8c77_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_8c77_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_8c77_return_output);

-- rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_cond,
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_iftrue,
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_iffalse,
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_8777
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_8777 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_8777_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_8777_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_8777_return_output);

-- rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_cond,
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_iftrue,
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_iffalse,
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_493d
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_493d : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_493d_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_493d_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_493d_return_output);

-- rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_cond,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_iftrue,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_iffalse,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_6132
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_6132 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_6132_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_6132_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_6132_return_output);

-- rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_cond,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_iftrue,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_iffalse,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_cc1e
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_cc1e : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_cc1e_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_cc1e_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_cc1e_return_output);

-- rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_cond,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_iftrue,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_iffalse,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_9d6a
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_9d6a : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_9d6a_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_9d6a_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_9d6a_return_output);

-- rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_cond,
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_iftrue,
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_iffalse,
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_8a43
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_8a43 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_8a43_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_8a43_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_8a43_return_output);

-- rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_cond,
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_iftrue,
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_iffalse,
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_814e
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_814e : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_814e_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_814e_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_814e_return_output);

-- rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_cond,
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_iftrue,
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_iffalse,
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_84b5
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_84b5 : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_84b5_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_84b5_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_84b5_return_output);

-- rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_cond,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_iftrue,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_iffalse,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_577e
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_577e : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_577e_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_577e_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_577e_return_output);

-- rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_cond,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_iftrue,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_iffalse,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_05b3
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_05b3 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_05b3_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_05b3_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_05b3_return_output);

-- rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_cond,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_iftrue,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_iffalse,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_a903
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_a903 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_a903_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_a903_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_a903_return_output);

-- rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_cond,
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_iftrue,
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_iffalse,
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_848c
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_848c : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_848c_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_848c_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_848c_return_output);

-- rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_cond,
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_iftrue,
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_iffalse,
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 elem_val,
 ref_toks_0,
 var_dim_0,
 -- All submodule outputs
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d584_return_output,
 rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_492e_return_output,
 rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_3a2b_return_output,
 rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_8c77_return_output,
 rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_8777_return_output,
 rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_493d_return_output,
 rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_6132_return_output,
 rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_cc1e_return_output,
 rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_9d6a_return_output,
 rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_8a43_return_output,
 rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_814e_return_output,
 rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_84b5_return_output,
 rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_577e_return_output,
 rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_05b3_return_output,
 rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_a903_return_output,
 rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_848c_return_output,
 rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_elem_val : unsigned(7 downto 0);
 variable VAR_ref_toks_0 : uint8_t_16;
 variable VAR_var_dim_0 : unsigned(3 downto 0);
 variable VAR_return_output : uint8_t_array_16_t;
 variable VAR_base : uint8_t_16;
 variable VAR_rv : uint8_t_array_16_t;
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l15_c15_3d3a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_8_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l16_c15_48ba_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l17_c15_117f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_11_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l18_c16_9d33_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_14_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l19_c16_7351_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l20_c15_3166_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l21_c15_752e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l22_c15_5c41_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_9_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l23_c15_6338_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_15_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l24_c16_4f26_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_12_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l25_c16_4933_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l26_c15_5f07_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l27_c15_f5ba_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l28_c15_72a0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_13_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l29_c16_a3b0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_10_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l30_c16_955f_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d584_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d584_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d584_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_492e_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_492e_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_492e_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_3a2b_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_3a2b_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_3a2b_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_8c77_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_8c77_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_8c77_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_8777_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_8777_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_8777_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_493d_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_493d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_493d_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_6132_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_6132_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_6132_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_cc1e_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_cc1e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_cc1e_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_9d6a_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_9d6a_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_9d6a_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_8a43_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_8a43_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_8a43_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_814e_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_814e_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_814e_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_84b5_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_84b5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_84b5_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_577e_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_577e_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_577e_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_05b3_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_05b3_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_05b3_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_a903_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_a903_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_a903_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_848c_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_848c_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_848c_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_eae2_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l129_c10_e0ef_return_output : uint8_t_array_16_t;
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_8c77_right := to_unsigned(11, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_814e_right := to_unsigned(12, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_848c_right := to_unsigned(10, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_3a2b_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_05b3_right := to_unsigned(7, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_493d_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_9d6a_right := to_unsigned(9, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_84b5_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_8a43_right := to_unsigned(15, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_cc1e_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_577e_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_a903_right := to_unsigned(13, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_6132_right := to_unsigned(6, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_492e_right := to_unsigned(8, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d584_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_8777_right := to_unsigned(14, 4);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_elem_val := elem_val;
     VAR_ref_toks_0 := ref_toks_0;
     VAR_var_dim_0 := var_dim_0;

     -- Submodule level 0
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_iftrue := VAR_elem_val;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_iftrue := VAR_elem_val;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_iftrue := VAR_elem_val;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_iftrue := VAR_elem_val;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_iftrue := VAR_elem_val;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_iftrue := VAR_elem_val;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_iftrue := VAR_elem_val;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_iftrue := VAR_elem_val;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_iftrue := VAR_elem_val;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_iftrue := VAR_elem_val;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_iftrue := VAR_elem_val;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_iftrue := VAR_elem_val;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_iftrue := VAR_elem_val;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_iftrue := VAR_elem_val;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_iftrue := VAR_elem_val;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_iftrue := VAR_elem_val;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_577e_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_05b3_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_a903_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_848c_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d584_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_492e_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_3a2b_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_8c77_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_8777_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_493d_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_6132_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_cc1e_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_9d6a_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_8a43_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_814e_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_84b5_left := VAR_var_dim_0;
     -- CONST_REF_RD_uint8_t_uint8_t_16_8_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l16_c15_48ba] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_8_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l16_c15_48ba_return_output := VAR_ref_toks_0(8);

     -- CONST_REF_RD_uint8_t_uint8_t_16_11_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l18_c16_9d33] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_11_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l18_c16_9d33_return_output := VAR_ref_toks_0(11);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_9d6a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_9d6a_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_9d6a_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_9d6a_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_9d6a_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_9d6a_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_9d6a_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_84b5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_84b5_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_84b5_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_84b5_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_84b5_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_84b5_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_84b5_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_6_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l21_c15_752e] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l21_c15_752e_return_output := VAR_ref_toks_0(6);

     -- CONST_REF_RD_uint8_t_uint8_t_16_2_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l15_c15_3d3a] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l15_c15_3d3a_return_output := VAR_ref_toks_0(2);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_cc1e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_cc1e_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_cc1e_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_cc1e_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_cc1e_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_cc1e_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_cc1e_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_5_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l17_c15_117f] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l17_c15_117f_return_output := VAR_ref_toks_0(5);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_a903] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_a903_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_a903_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_a903_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_a903_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_a903_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_a903_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_6132] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_6132_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_6132_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_6132_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_6132_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_6132_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_6132_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_3_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l22_c15_5c41] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l22_c15_5c41_return_output := VAR_ref_toks_0(3);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_814e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_814e_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_814e_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_814e_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_814e_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_814e_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_814e_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_15_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l24_c16_4f26] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_15_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l24_c16_4f26_return_output := VAR_ref_toks_0(15);

     -- CONST_REF_RD_uint8_t_uint8_t_16_13_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l29_c16_a3b0] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_13_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l29_c16_a3b0_return_output := VAR_ref_toks_0(13);

     -- CONST_REF_RD_uint8_t_uint8_t_16_14_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l19_c16_7351] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_14_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l19_c16_7351_return_output := VAR_ref_toks_0(14);

     -- CONST_REF_RD_uint8_t_uint8_t_16_4_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l27_c15_f5ba] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l27_c15_f5ba_return_output := VAR_ref_toks_0(4);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d584] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d584_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d584_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d584_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d584_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d584_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d584_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_8a43] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_8a43_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_8a43_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_8a43_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_8a43_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_8a43_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_8a43_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_0_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l20_c15_3166] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l20_c15_3166_return_output := VAR_ref_toks_0(0);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_05b3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_05b3_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_05b3_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_05b3_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_05b3_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_05b3_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_05b3_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_492e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_492e_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_492e_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_492e_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_492e_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_492e_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_492e_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_8c77] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_8c77_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_8c77_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_8c77_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_8c77_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_8c77_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_8c77_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_3a2b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_3a2b_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_3a2b_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_3a2b_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_3a2b_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_3a2b_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_3a2b_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_1_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l26_c15_5f07] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l26_c15_5f07_return_output := VAR_ref_toks_0(1);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_493d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_493d_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_493d_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_493d_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_493d_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_493d_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_493d_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_577e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_577e_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_577e_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_577e_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_577e_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_577e_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_577e_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_848c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_848c_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_848c_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_848c_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_848c_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_848c_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_848c_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_9_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l23_c15_6338] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_9_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l23_c15_6338_return_output := VAR_ref_toks_0(9);

     -- CONST_REF_RD_uint8_t_uint8_t_16_7_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l28_c15_72a0] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l28_c15_72a0_return_output := VAR_ref_toks_0(7);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_8777] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_8777_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_8777_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_8777_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_8777_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_8777_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_8777_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_12_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l25_c16_4933] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_12_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l25_c16_4933_return_output := VAR_ref_toks_0(12);

     -- CONST_REF_RD_uint8_t_uint8_t_16_10_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l30_c16_955f] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_10_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l30_c16_955f_return_output := VAR_ref_toks_0(10);

     -- Submodule level 1
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_577e_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_05b3_return_output;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_a903_return_output;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_848c_return_output;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_d584_return_output;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_492e_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_3a2b_return_output;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_8c77_return_output;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_8777_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_493d_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_6132_return_output;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_cc1e_return_output;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_9d6a_return_output;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_8a43_return_output;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_814e_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_84b5_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l20_c15_3166_return_output;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_10_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l30_c16_955f_return_output;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_11_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l18_c16_9d33_return_output;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_12_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l25_c16_4933_return_output;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_13_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l29_c16_a3b0_return_output;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_14_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l19_c16_7351_return_output;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_15_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l24_c16_4f26_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l26_c15_5f07_return_output;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l15_c15_3d3a_return_output;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l22_c15_5c41_return_output;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l27_c15_f5ba_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l17_c15_117f_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l21_c15_752e_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l28_c15_72a0_return_output;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_8_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l16_c15_48ba_return_output;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_9_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l23_c15_6338_return_output;
     -- rv_data_10_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf] LATENCY=0
     -- Inputs
     rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_cond <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_cond;
     rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_iftrue <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_iftrue;
     rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_iffalse <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_iffalse;
     -- Outputs
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_return_output := rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_return_output;

     -- rv_data_4_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741] LATENCY=0
     -- Inputs
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_cond <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_cond;
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_iftrue <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_iftrue;
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_iffalse <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_iffalse;
     -- Outputs
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_return_output := rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_return_output;

     -- rv_data_6_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506] LATENCY=0
     -- Inputs
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_cond <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_cond;
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_iftrue <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_iftrue;
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_iffalse <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_iffalse;
     -- Outputs
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_return_output := rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_return_output;

     -- rv_data_13_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b] LATENCY=0
     -- Inputs
     rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_cond <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_cond;
     rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_iftrue <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_iftrue;
     rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_iffalse <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_iffalse;
     -- Outputs
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_return_output := rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_return_output;

     -- rv_data_14_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431] LATENCY=0
     -- Inputs
     rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_cond <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_cond;
     rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_iftrue <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_iftrue;
     rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_iffalse <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_iffalse;
     -- Outputs
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_return_output := rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_return_output;

     -- rv_data_12_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3] LATENCY=0
     -- Inputs
     rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_cond <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_cond;
     rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_iftrue <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_iftrue;
     rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_iffalse <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_iffalse;
     -- Outputs
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_return_output := rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_return_output;

     -- rv_data_0_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c] LATENCY=0
     -- Inputs
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_cond <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_cond;
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_iftrue <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_iftrue;
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_iffalse <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_iffalse;
     -- Outputs
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_return_output := rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_return_output;

     -- rv_data_3_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8] LATENCY=0
     -- Inputs
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_cond <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_cond;
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_iftrue <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_iftrue;
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_iffalse <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_iffalse;
     -- Outputs
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_return_output := rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_return_output;

     -- rv_data_11_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171] LATENCY=0
     -- Inputs
     rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_cond <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_cond;
     rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_iftrue <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_iftrue;
     rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_iffalse <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_iffalse;
     -- Outputs
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_return_output := rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_return_output;

     -- rv_data_7_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778] LATENCY=0
     -- Inputs
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_cond <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_cond;
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_iftrue <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_iftrue;
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_iffalse <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_iffalse;
     -- Outputs
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_return_output := rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_return_output;

     -- rv_data_1_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d] LATENCY=0
     -- Inputs
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_cond <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_cond;
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_iftrue <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_iftrue;
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_iffalse <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_iffalse;
     -- Outputs
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_return_output := rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_return_output;

     -- rv_data_15_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c] LATENCY=0
     -- Inputs
     rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_cond <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_cond;
     rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_iftrue <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_iftrue;
     rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_iffalse <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_iffalse;
     -- Outputs
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_return_output := rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_return_output;

     -- rv_data_2_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a] LATENCY=0
     -- Inputs
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_cond <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_cond;
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_iftrue <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_iftrue;
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_iffalse <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_iffalse;
     -- Outputs
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_return_output := rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_return_output;

     -- rv_data_5_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43] LATENCY=0
     -- Inputs
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_cond <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_cond;
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_iftrue <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_iftrue;
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_iffalse <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_iffalse;
     -- Outputs
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_return_output := rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_return_output;

     -- rv_data_8_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d] LATENCY=0
     -- Inputs
     rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_cond <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_cond;
     rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_iftrue <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_iftrue;
     rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_iffalse <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_iffalse;
     -- Outputs
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_return_output := rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_return_output;

     -- rv_data_9_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea] LATENCY=0
     -- Inputs
     rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_cond <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_cond;
     rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_iftrue <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_iftrue;
     rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_iffalse <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_iffalse;
     -- Outputs
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_return_output := rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_return_output;

     -- Submodule level 2
     -- CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_eae2[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l129_c10_e0ef] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_eae2_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l129_c10_e0ef_return_output := CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_eae2(
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_2c8a_return_output,
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4f6d_return_output,
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_0a43_return_output,
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_e171_return_output,
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_5431_return_output,
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_589c_return_output,
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_1506_return_output,
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_67d8_return_output,
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_67ea_return_output,
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_920c_return_output,
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_b0c3_return_output,
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_995d_return_output,
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_6741_return_output,
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_d778_return_output,
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_c35b_return_output,
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_48cf_return_output);

     -- Submodule level 3
     VAR_return_output := VAR_CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_eae2_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l129_c10_e0ef_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
