-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 134
entity uint8_mux128_0CLK_9347d63d is
port(
 sel : in unsigned(6 downto 0);
 in0 : in unsigned(7 downto 0);
 in1 : in unsigned(7 downto 0);
 in2 : in unsigned(7 downto 0);
 in3 : in unsigned(7 downto 0);
 in4 : in unsigned(7 downto 0);
 in5 : in unsigned(7 downto 0);
 in6 : in unsigned(7 downto 0);
 in7 : in unsigned(7 downto 0);
 in8 : in unsigned(7 downto 0);
 in9 : in unsigned(7 downto 0);
 in10 : in unsigned(7 downto 0);
 in11 : in unsigned(7 downto 0);
 in12 : in unsigned(7 downto 0);
 in13 : in unsigned(7 downto 0);
 in14 : in unsigned(7 downto 0);
 in15 : in unsigned(7 downto 0);
 in16 : in unsigned(7 downto 0);
 in17 : in unsigned(7 downto 0);
 in18 : in unsigned(7 downto 0);
 in19 : in unsigned(7 downto 0);
 in20 : in unsigned(7 downto 0);
 in21 : in unsigned(7 downto 0);
 in22 : in unsigned(7 downto 0);
 in23 : in unsigned(7 downto 0);
 in24 : in unsigned(7 downto 0);
 in25 : in unsigned(7 downto 0);
 in26 : in unsigned(7 downto 0);
 in27 : in unsigned(7 downto 0);
 in28 : in unsigned(7 downto 0);
 in29 : in unsigned(7 downto 0);
 in30 : in unsigned(7 downto 0);
 in31 : in unsigned(7 downto 0);
 in32 : in unsigned(7 downto 0);
 in33 : in unsigned(7 downto 0);
 in34 : in unsigned(7 downto 0);
 in35 : in unsigned(7 downto 0);
 in36 : in unsigned(7 downto 0);
 in37 : in unsigned(7 downto 0);
 in38 : in unsigned(7 downto 0);
 in39 : in unsigned(7 downto 0);
 in40 : in unsigned(7 downto 0);
 in41 : in unsigned(7 downto 0);
 in42 : in unsigned(7 downto 0);
 in43 : in unsigned(7 downto 0);
 in44 : in unsigned(7 downto 0);
 in45 : in unsigned(7 downto 0);
 in46 : in unsigned(7 downto 0);
 in47 : in unsigned(7 downto 0);
 in48 : in unsigned(7 downto 0);
 in49 : in unsigned(7 downto 0);
 in50 : in unsigned(7 downto 0);
 in51 : in unsigned(7 downto 0);
 in52 : in unsigned(7 downto 0);
 in53 : in unsigned(7 downto 0);
 in54 : in unsigned(7 downto 0);
 in55 : in unsigned(7 downto 0);
 in56 : in unsigned(7 downto 0);
 in57 : in unsigned(7 downto 0);
 in58 : in unsigned(7 downto 0);
 in59 : in unsigned(7 downto 0);
 in60 : in unsigned(7 downto 0);
 in61 : in unsigned(7 downto 0);
 in62 : in unsigned(7 downto 0);
 in63 : in unsigned(7 downto 0);
 in64 : in unsigned(7 downto 0);
 in65 : in unsigned(7 downto 0);
 in66 : in unsigned(7 downto 0);
 in67 : in unsigned(7 downto 0);
 in68 : in unsigned(7 downto 0);
 in69 : in unsigned(7 downto 0);
 in70 : in unsigned(7 downto 0);
 in71 : in unsigned(7 downto 0);
 in72 : in unsigned(7 downto 0);
 in73 : in unsigned(7 downto 0);
 in74 : in unsigned(7 downto 0);
 in75 : in unsigned(7 downto 0);
 in76 : in unsigned(7 downto 0);
 in77 : in unsigned(7 downto 0);
 in78 : in unsigned(7 downto 0);
 in79 : in unsigned(7 downto 0);
 in80 : in unsigned(7 downto 0);
 in81 : in unsigned(7 downto 0);
 in82 : in unsigned(7 downto 0);
 in83 : in unsigned(7 downto 0);
 in84 : in unsigned(7 downto 0);
 in85 : in unsigned(7 downto 0);
 in86 : in unsigned(7 downto 0);
 in87 : in unsigned(7 downto 0);
 in88 : in unsigned(7 downto 0);
 in89 : in unsigned(7 downto 0);
 in90 : in unsigned(7 downto 0);
 in91 : in unsigned(7 downto 0);
 in92 : in unsigned(7 downto 0);
 in93 : in unsigned(7 downto 0);
 in94 : in unsigned(7 downto 0);
 in95 : in unsigned(7 downto 0);
 in96 : in unsigned(7 downto 0);
 in97 : in unsigned(7 downto 0);
 in98 : in unsigned(7 downto 0);
 in99 : in unsigned(7 downto 0);
 in100 : in unsigned(7 downto 0);
 in101 : in unsigned(7 downto 0);
 in102 : in unsigned(7 downto 0);
 in103 : in unsigned(7 downto 0);
 in104 : in unsigned(7 downto 0);
 in105 : in unsigned(7 downto 0);
 in106 : in unsigned(7 downto 0);
 in107 : in unsigned(7 downto 0);
 in108 : in unsigned(7 downto 0);
 in109 : in unsigned(7 downto 0);
 in110 : in unsigned(7 downto 0);
 in111 : in unsigned(7 downto 0);
 in112 : in unsigned(7 downto 0);
 in113 : in unsigned(7 downto 0);
 in114 : in unsigned(7 downto 0);
 in115 : in unsigned(7 downto 0);
 in116 : in unsigned(7 downto 0);
 in117 : in unsigned(7 downto 0);
 in118 : in unsigned(7 downto 0);
 in119 : in unsigned(7 downto 0);
 in120 : in unsigned(7 downto 0);
 in121 : in unsigned(7 downto 0);
 in122 : in unsigned(7 downto 0);
 in123 : in unsigned(7 downto 0);
 in124 : in unsigned(7 downto 0);
 in125 : in unsigned(7 downto 0);
 in126 : in unsigned(7 downto 0);
 in127 : in unsigned(7 downto 0);
 return_output : out unsigned(7 downto 0));
end uint8_mux128_0CLK_9347d63d;
architecture arch of uint8_mux128_0CLK_9347d63d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- layer0_node0_MUX[bit_math_h_l18_c3_ce9b]
signal layer0_node0_MUX_bit_math_h_l18_c3_ce9b_cond : unsigned(0 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_ce9b_iftrue : unsigned(7 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_ce9b_iffalse : unsigned(7 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_ce9b_return_output : unsigned(7 downto 0);

-- layer0_node1_MUX[bit_math_h_l29_c3_0e94]
signal layer0_node1_MUX_bit_math_h_l29_c3_0e94_cond : unsigned(0 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_0e94_iftrue : unsigned(7 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_0e94_iffalse : unsigned(7 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_0e94_return_output : unsigned(7 downto 0);

-- layer0_node2_MUX[bit_math_h_l40_c3_e2d9]
signal layer0_node2_MUX_bit_math_h_l40_c3_e2d9_cond : unsigned(0 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_e2d9_iftrue : unsigned(7 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_e2d9_iffalse : unsigned(7 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_e2d9_return_output : unsigned(7 downto 0);

-- layer0_node3_MUX[bit_math_h_l51_c3_edc9]
signal layer0_node3_MUX_bit_math_h_l51_c3_edc9_cond : unsigned(0 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_edc9_iftrue : unsigned(7 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_edc9_iffalse : unsigned(7 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_edc9_return_output : unsigned(7 downto 0);

-- layer0_node4_MUX[bit_math_h_l62_c3_f389]
signal layer0_node4_MUX_bit_math_h_l62_c3_f389_cond : unsigned(0 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_f389_iftrue : unsigned(7 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_f389_iffalse : unsigned(7 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_f389_return_output : unsigned(7 downto 0);

-- layer0_node5_MUX[bit_math_h_l73_c3_d655]
signal layer0_node5_MUX_bit_math_h_l73_c3_d655_cond : unsigned(0 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_d655_iftrue : unsigned(7 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_d655_iffalse : unsigned(7 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_d655_return_output : unsigned(7 downto 0);

-- layer0_node6_MUX[bit_math_h_l84_c3_5cd3]
signal layer0_node6_MUX_bit_math_h_l84_c3_5cd3_cond : unsigned(0 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_5cd3_iftrue : unsigned(7 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_5cd3_iffalse : unsigned(7 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_5cd3_return_output : unsigned(7 downto 0);

-- layer0_node7_MUX[bit_math_h_l95_c3_5030]
signal layer0_node7_MUX_bit_math_h_l95_c3_5030_cond : unsigned(0 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_5030_iftrue : unsigned(7 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_5030_iffalse : unsigned(7 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_5030_return_output : unsigned(7 downto 0);

-- layer0_node8_MUX[bit_math_h_l106_c3_32cb]
signal layer0_node8_MUX_bit_math_h_l106_c3_32cb_cond : unsigned(0 downto 0);
signal layer0_node8_MUX_bit_math_h_l106_c3_32cb_iftrue : unsigned(7 downto 0);
signal layer0_node8_MUX_bit_math_h_l106_c3_32cb_iffalse : unsigned(7 downto 0);
signal layer0_node8_MUX_bit_math_h_l106_c3_32cb_return_output : unsigned(7 downto 0);

-- layer0_node9_MUX[bit_math_h_l117_c3_4b42]
signal layer0_node9_MUX_bit_math_h_l117_c3_4b42_cond : unsigned(0 downto 0);
signal layer0_node9_MUX_bit_math_h_l117_c3_4b42_iftrue : unsigned(7 downto 0);
signal layer0_node9_MUX_bit_math_h_l117_c3_4b42_iffalse : unsigned(7 downto 0);
signal layer0_node9_MUX_bit_math_h_l117_c3_4b42_return_output : unsigned(7 downto 0);

-- layer0_node10_MUX[bit_math_h_l128_c3_06f3]
signal layer0_node10_MUX_bit_math_h_l128_c3_06f3_cond : unsigned(0 downto 0);
signal layer0_node10_MUX_bit_math_h_l128_c3_06f3_iftrue : unsigned(7 downto 0);
signal layer0_node10_MUX_bit_math_h_l128_c3_06f3_iffalse : unsigned(7 downto 0);
signal layer0_node10_MUX_bit_math_h_l128_c3_06f3_return_output : unsigned(7 downto 0);

-- layer0_node11_MUX[bit_math_h_l139_c3_dbfc]
signal layer0_node11_MUX_bit_math_h_l139_c3_dbfc_cond : unsigned(0 downto 0);
signal layer0_node11_MUX_bit_math_h_l139_c3_dbfc_iftrue : unsigned(7 downto 0);
signal layer0_node11_MUX_bit_math_h_l139_c3_dbfc_iffalse : unsigned(7 downto 0);
signal layer0_node11_MUX_bit_math_h_l139_c3_dbfc_return_output : unsigned(7 downto 0);

-- layer0_node12_MUX[bit_math_h_l150_c3_6613]
signal layer0_node12_MUX_bit_math_h_l150_c3_6613_cond : unsigned(0 downto 0);
signal layer0_node12_MUX_bit_math_h_l150_c3_6613_iftrue : unsigned(7 downto 0);
signal layer0_node12_MUX_bit_math_h_l150_c3_6613_iffalse : unsigned(7 downto 0);
signal layer0_node12_MUX_bit_math_h_l150_c3_6613_return_output : unsigned(7 downto 0);

-- layer0_node13_MUX[bit_math_h_l161_c3_fd42]
signal layer0_node13_MUX_bit_math_h_l161_c3_fd42_cond : unsigned(0 downto 0);
signal layer0_node13_MUX_bit_math_h_l161_c3_fd42_iftrue : unsigned(7 downto 0);
signal layer0_node13_MUX_bit_math_h_l161_c3_fd42_iffalse : unsigned(7 downto 0);
signal layer0_node13_MUX_bit_math_h_l161_c3_fd42_return_output : unsigned(7 downto 0);

-- layer0_node14_MUX[bit_math_h_l172_c3_154a]
signal layer0_node14_MUX_bit_math_h_l172_c3_154a_cond : unsigned(0 downto 0);
signal layer0_node14_MUX_bit_math_h_l172_c3_154a_iftrue : unsigned(7 downto 0);
signal layer0_node14_MUX_bit_math_h_l172_c3_154a_iffalse : unsigned(7 downto 0);
signal layer0_node14_MUX_bit_math_h_l172_c3_154a_return_output : unsigned(7 downto 0);

-- layer0_node15_MUX[bit_math_h_l183_c3_5274]
signal layer0_node15_MUX_bit_math_h_l183_c3_5274_cond : unsigned(0 downto 0);
signal layer0_node15_MUX_bit_math_h_l183_c3_5274_iftrue : unsigned(7 downto 0);
signal layer0_node15_MUX_bit_math_h_l183_c3_5274_iffalse : unsigned(7 downto 0);
signal layer0_node15_MUX_bit_math_h_l183_c3_5274_return_output : unsigned(7 downto 0);

-- layer0_node16_MUX[bit_math_h_l194_c3_7a7d]
signal layer0_node16_MUX_bit_math_h_l194_c3_7a7d_cond : unsigned(0 downto 0);
signal layer0_node16_MUX_bit_math_h_l194_c3_7a7d_iftrue : unsigned(7 downto 0);
signal layer0_node16_MUX_bit_math_h_l194_c3_7a7d_iffalse : unsigned(7 downto 0);
signal layer0_node16_MUX_bit_math_h_l194_c3_7a7d_return_output : unsigned(7 downto 0);

-- layer0_node17_MUX[bit_math_h_l205_c3_42ac]
signal layer0_node17_MUX_bit_math_h_l205_c3_42ac_cond : unsigned(0 downto 0);
signal layer0_node17_MUX_bit_math_h_l205_c3_42ac_iftrue : unsigned(7 downto 0);
signal layer0_node17_MUX_bit_math_h_l205_c3_42ac_iffalse : unsigned(7 downto 0);
signal layer0_node17_MUX_bit_math_h_l205_c3_42ac_return_output : unsigned(7 downto 0);

-- layer0_node18_MUX[bit_math_h_l216_c3_b8f1]
signal layer0_node18_MUX_bit_math_h_l216_c3_b8f1_cond : unsigned(0 downto 0);
signal layer0_node18_MUX_bit_math_h_l216_c3_b8f1_iftrue : unsigned(7 downto 0);
signal layer0_node18_MUX_bit_math_h_l216_c3_b8f1_iffalse : unsigned(7 downto 0);
signal layer0_node18_MUX_bit_math_h_l216_c3_b8f1_return_output : unsigned(7 downto 0);

-- layer0_node19_MUX[bit_math_h_l227_c3_0b12]
signal layer0_node19_MUX_bit_math_h_l227_c3_0b12_cond : unsigned(0 downto 0);
signal layer0_node19_MUX_bit_math_h_l227_c3_0b12_iftrue : unsigned(7 downto 0);
signal layer0_node19_MUX_bit_math_h_l227_c3_0b12_iffalse : unsigned(7 downto 0);
signal layer0_node19_MUX_bit_math_h_l227_c3_0b12_return_output : unsigned(7 downto 0);

-- layer0_node20_MUX[bit_math_h_l238_c3_091e]
signal layer0_node20_MUX_bit_math_h_l238_c3_091e_cond : unsigned(0 downto 0);
signal layer0_node20_MUX_bit_math_h_l238_c3_091e_iftrue : unsigned(7 downto 0);
signal layer0_node20_MUX_bit_math_h_l238_c3_091e_iffalse : unsigned(7 downto 0);
signal layer0_node20_MUX_bit_math_h_l238_c3_091e_return_output : unsigned(7 downto 0);

-- layer0_node21_MUX[bit_math_h_l249_c3_44d2]
signal layer0_node21_MUX_bit_math_h_l249_c3_44d2_cond : unsigned(0 downto 0);
signal layer0_node21_MUX_bit_math_h_l249_c3_44d2_iftrue : unsigned(7 downto 0);
signal layer0_node21_MUX_bit_math_h_l249_c3_44d2_iffalse : unsigned(7 downto 0);
signal layer0_node21_MUX_bit_math_h_l249_c3_44d2_return_output : unsigned(7 downto 0);

-- layer0_node22_MUX[bit_math_h_l260_c3_db28]
signal layer0_node22_MUX_bit_math_h_l260_c3_db28_cond : unsigned(0 downto 0);
signal layer0_node22_MUX_bit_math_h_l260_c3_db28_iftrue : unsigned(7 downto 0);
signal layer0_node22_MUX_bit_math_h_l260_c3_db28_iffalse : unsigned(7 downto 0);
signal layer0_node22_MUX_bit_math_h_l260_c3_db28_return_output : unsigned(7 downto 0);

-- layer0_node23_MUX[bit_math_h_l271_c3_0038]
signal layer0_node23_MUX_bit_math_h_l271_c3_0038_cond : unsigned(0 downto 0);
signal layer0_node23_MUX_bit_math_h_l271_c3_0038_iftrue : unsigned(7 downto 0);
signal layer0_node23_MUX_bit_math_h_l271_c3_0038_iffalse : unsigned(7 downto 0);
signal layer0_node23_MUX_bit_math_h_l271_c3_0038_return_output : unsigned(7 downto 0);

-- layer0_node24_MUX[bit_math_h_l282_c3_1d56]
signal layer0_node24_MUX_bit_math_h_l282_c3_1d56_cond : unsigned(0 downto 0);
signal layer0_node24_MUX_bit_math_h_l282_c3_1d56_iftrue : unsigned(7 downto 0);
signal layer0_node24_MUX_bit_math_h_l282_c3_1d56_iffalse : unsigned(7 downto 0);
signal layer0_node24_MUX_bit_math_h_l282_c3_1d56_return_output : unsigned(7 downto 0);

-- layer0_node25_MUX[bit_math_h_l293_c3_fa3c]
signal layer0_node25_MUX_bit_math_h_l293_c3_fa3c_cond : unsigned(0 downto 0);
signal layer0_node25_MUX_bit_math_h_l293_c3_fa3c_iftrue : unsigned(7 downto 0);
signal layer0_node25_MUX_bit_math_h_l293_c3_fa3c_iffalse : unsigned(7 downto 0);
signal layer0_node25_MUX_bit_math_h_l293_c3_fa3c_return_output : unsigned(7 downto 0);

-- layer0_node26_MUX[bit_math_h_l304_c3_220e]
signal layer0_node26_MUX_bit_math_h_l304_c3_220e_cond : unsigned(0 downto 0);
signal layer0_node26_MUX_bit_math_h_l304_c3_220e_iftrue : unsigned(7 downto 0);
signal layer0_node26_MUX_bit_math_h_l304_c3_220e_iffalse : unsigned(7 downto 0);
signal layer0_node26_MUX_bit_math_h_l304_c3_220e_return_output : unsigned(7 downto 0);

-- layer0_node27_MUX[bit_math_h_l315_c3_37d2]
signal layer0_node27_MUX_bit_math_h_l315_c3_37d2_cond : unsigned(0 downto 0);
signal layer0_node27_MUX_bit_math_h_l315_c3_37d2_iftrue : unsigned(7 downto 0);
signal layer0_node27_MUX_bit_math_h_l315_c3_37d2_iffalse : unsigned(7 downto 0);
signal layer0_node27_MUX_bit_math_h_l315_c3_37d2_return_output : unsigned(7 downto 0);

-- layer0_node28_MUX[bit_math_h_l326_c3_af14]
signal layer0_node28_MUX_bit_math_h_l326_c3_af14_cond : unsigned(0 downto 0);
signal layer0_node28_MUX_bit_math_h_l326_c3_af14_iftrue : unsigned(7 downto 0);
signal layer0_node28_MUX_bit_math_h_l326_c3_af14_iffalse : unsigned(7 downto 0);
signal layer0_node28_MUX_bit_math_h_l326_c3_af14_return_output : unsigned(7 downto 0);

-- layer0_node29_MUX[bit_math_h_l337_c3_d491]
signal layer0_node29_MUX_bit_math_h_l337_c3_d491_cond : unsigned(0 downto 0);
signal layer0_node29_MUX_bit_math_h_l337_c3_d491_iftrue : unsigned(7 downto 0);
signal layer0_node29_MUX_bit_math_h_l337_c3_d491_iffalse : unsigned(7 downto 0);
signal layer0_node29_MUX_bit_math_h_l337_c3_d491_return_output : unsigned(7 downto 0);

-- layer0_node30_MUX[bit_math_h_l348_c3_46cf]
signal layer0_node30_MUX_bit_math_h_l348_c3_46cf_cond : unsigned(0 downto 0);
signal layer0_node30_MUX_bit_math_h_l348_c3_46cf_iftrue : unsigned(7 downto 0);
signal layer0_node30_MUX_bit_math_h_l348_c3_46cf_iffalse : unsigned(7 downto 0);
signal layer0_node30_MUX_bit_math_h_l348_c3_46cf_return_output : unsigned(7 downto 0);

-- layer0_node31_MUX[bit_math_h_l359_c3_1ee6]
signal layer0_node31_MUX_bit_math_h_l359_c3_1ee6_cond : unsigned(0 downto 0);
signal layer0_node31_MUX_bit_math_h_l359_c3_1ee6_iftrue : unsigned(7 downto 0);
signal layer0_node31_MUX_bit_math_h_l359_c3_1ee6_iffalse : unsigned(7 downto 0);
signal layer0_node31_MUX_bit_math_h_l359_c3_1ee6_return_output : unsigned(7 downto 0);

-- layer0_node32_MUX[bit_math_h_l370_c3_ee39]
signal layer0_node32_MUX_bit_math_h_l370_c3_ee39_cond : unsigned(0 downto 0);
signal layer0_node32_MUX_bit_math_h_l370_c3_ee39_iftrue : unsigned(7 downto 0);
signal layer0_node32_MUX_bit_math_h_l370_c3_ee39_iffalse : unsigned(7 downto 0);
signal layer0_node32_MUX_bit_math_h_l370_c3_ee39_return_output : unsigned(7 downto 0);

-- layer0_node33_MUX[bit_math_h_l381_c3_f57d]
signal layer0_node33_MUX_bit_math_h_l381_c3_f57d_cond : unsigned(0 downto 0);
signal layer0_node33_MUX_bit_math_h_l381_c3_f57d_iftrue : unsigned(7 downto 0);
signal layer0_node33_MUX_bit_math_h_l381_c3_f57d_iffalse : unsigned(7 downto 0);
signal layer0_node33_MUX_bit_math_h_l381_c3_f57d_return_output : unsigned(7 downto 0);

-- layer0_node34_MUX[bit_math_h_l392_c3_8d4e]
signal layer0_node34_MUX_bit_math_h_l392_c3_8d4e_cond : unsigned(0 downto 0);
signal layer0_node34_MUX_bit_math_h_l392_c3_8d4e_iftrue : unsigned(7 downto 0);
signal layer0_node34_MUX_bit_math_h_l392_c3_8d4e_iffalse : unsigned(7 downto 0);
signal layer0_node34_MUX_bit_math_h_l392_c3_8d4e_return_output : unsigned(7 downto 0);

-- layer0_node35_MUX[bit_math_h_l403_c3_fa1f]
signal layer0_node35_MUX_bit_math_h_l403_c3_fa1f_cond : unsigned(0 downto 0);
signal layer0_node35_MUX_bit_math_h_l403_c3_fa1f_iftrue : unsigned(7 downto 0);
signal layer0_node35_MUX_bit_math_h_l403_c3_fa1f_iffalse : unsigned(7 downto 0);
signal layer0_node35_MUX_bit_math_h_l403_c3_fa1f_return_output : unsigned(7 downto 0);

-- layer0_node36_MUX[bit_math_h_l414_c3_39b4]
signal layer0_node36_MUX_bit_math_h_l414_c3_39b4_cond : unsigned(0 downto 0);
signal layer0_node36_MUX_bit_math_h_l414_c3_39b4_iftrue : unsigned(7 downto 0);
signal layer0_node36_MUX_bit_math_h_l414_c3_39b4_iffalse : unsigned(7 downto 0);
signal layer0_node36_MUX_bit_math_h_l414_c3_39b4_return_output : unsigned(7 downto 0);

-- layer0_node37_MUX[bit_math_h_l425_c3_3900]
signal layer0_node37_MUX_bit_math_h_l425_c3_3900_cond : unsigned(0 downto 0);
signal layer0_node37_MUX_bit_math_h_l425_c3_3900_iftrue : unsigned(7 downto 0);
signal layer0_node37_MUX_bit_math_h_l425_c3_3900_iffalse : unsigned(7 downto 0);
signal layer0_node37_MUX_bit_math_h_l425_c3_3900_return_output : unsigned(7 downto 0);

-- layer0_node38_MUX[bit_math_h_l436_c3_bea2]
signal layer0_node38_MUX_bit_math_h_l436_c3_bea2_cond : unsigned(0 downto 0);
signal layer0_node38_MUX_bit_math_h_l436_c3_bea2_iftrue : unsigned(7 downto 0);
signal layer0_node38_MUX_bit_math_h_l436_c3_bea2_iffalse : unsigned(7 downto 0);
signal layer0_node38_MUX_bit_math_h_l436_c3_bea2_return_output : unsigned(7 downto 0);

-- layer0_node39_MUX[bit_math_h_l447_c3_3acc]
signal layer0_node39_MUX_bit_math_h_l447_c3_3acc_cond : unsigned(0 downto 0);
signal layer0_node39_MUX_bit_math_h_l447_c3_3acc_iftrue : unsigned(7 downto 0);
signal layer0_node39_MUX_bit_math_h_l447_c3_3acc_iffalse : unsigned(7 downto 0);
signal layer0_node39_MUX_bit_math_h_l447_c3_3acc_return_output : unsigned(7 downto 0);

-- layer0_node40_MUX[bit_math_h_l458_c3_f867]
signal layer0_node40_MUX_bit_math_h_l458_c3_f867_cond : unsigned(0 downto 0);
signal layer0_node40_MUX_bit_math_h_l458_c3_f867_iftrue : unsigned(7 downto 0);
signal layer0_node40_MUX_bit_math_h_l458_c3_f867_iffalse : unsigned(7 downto 0);
signal layer0_node40_MUX_bit_math_h_l458_c3_f867_return_output : unsigned(7 downto 0);

-- layer0_node41_MUX[bit_math_h_l469_c3_2ffe]
signal layer0_node41_MUX_bit_math_h_l469_c3_2ffe_cond : unsigned(0 downto 0);
signal layer0_node41_MUX_bit_math_h_l469_c3_2ffe_iftrue : unsigned(7 downto 0);
signal layer0_node41_MUX_bit_math_h_l469_c3_2ffe_iffalse : unsigned(7 downto 0);
signal layer0_node41_MUX_bit_math_h_l469_c3_2ffe_return_output : unsigned(7 downto 0);

-- layer0_node42_MUX[bit_math_h_l480_c3_1c62]
signal layer0_node42_MUX_bit_math_h_l480_c3_1c62_cond : unsigned(0 downto 0);
signal layer0_node42_MUX_bit_math_h_l480_c3_1c62_iftrue : unsigned(7 downto 0);
signal layer0_node42_MUX_bit_math_h_l480_c3_1c62_iffalse : unsigned(7 downto 0);
signal layer0_node42_MUX_bit_math_h_l480_c3_1c62_return_output : unsigned(7 downto 0);

-- layer0_node43_MUX[bit_math_h_l491_c3_7943]
signal layer0_node43_MUX_bit_math_h_l491_c3_7943_cond : unsigned(0 downto 0);
signal layer0_node43_MUX_bit_math_h_l491_c3_7943_iftrue : unsigned(7 downto 0);
signal layer0_node43_MUX_bit_math_h_l491_c3_7943_iffalse : unsigned(7 downto 0);
signal layer0_node43_MUX_bit_math_h_l491_c3_7943_return_output : unsigned(7 downto 0);

-- layer0_node44_MUX[bit_math_h_l502_c3_15dc]
signal layer0_node44_MUX_bit_math_h_l502_c3_15dc_cond : unsigned(0 downto 0);
signal layer0_node44_MUX_bit_math_h_l502_c3_15dc_iftrue : unsigned(7 downto 0);
signal layer0_node44_MUX_bit_math_h_l502_c3_15dc_iffalse : unsigned(7 downto 0);
signal layer0_node44_MUX_bit_math_h_l502_c3_15dc_return_output : unsigned(7 downto 0);

-- layer0_node45_MUX[bit_math_h_l513_c3_d638]
signal layer0_node45_MUX_bit_math_h_l513_c3_d638_cond : unsigned(0 downto 0);
signal layer0_node45_MUX_bit_math_h_l513_c3_d638_iftrue : unsigned(7 downto 0);
signal layer0_node45_MUX_bit_math_h_l513_c3_d638_iffalse : unsigned(7 downto 0);
signal layer0_node45_MUX_bit_math_h_l513_c3_d638_return_output : unsigned(7 downto 0);

-- layer0_node46_MUX[bit_math_h_l524_c3_fdc0]
signal layer0_node46_MUX_bit_math_h_l524_c3_fdc0_cond : unsigned(0 downto 0);
signal layer0_node46_MUX_bit_math_h_l524_c3_fdc0_iftrue : unsigned(7 downto 0);
signal layer0_node46_MUX_bit_math_h_l524_c3_fdc0_iffalse : unsigned(7 downto 0);
signal layer0_node46_MUX_bit_math_h_l524_c3_fdc0_return_output : unsigned(7 downto 0);

-- layer0_node47_MUX[bit_math_h_l535_c3_1640]
signal layer0_node47_MUX_bit_math_h_l535_c3_1640_cond : unsigned(0 downto 0);
signal layer0_node47_MUX_bit_math_h_l535_c3_1640_iftrue : unsigned(7 downto 0);
signal layer0_node47_MUX_bit_math_h_l535_c3_1640_iffalse : unsigned(7 downto 0);
signal layer0_node47_MUX_bit_math_h_l535_c3_1640_return_output : unsigned(7 downto 0);

-- layer0_node48_MUX[bit_math_h_l546_c3_b0f6]
signal layer0_node48_MUX_bit_math_h_l546_c3_b0f6_cond : unsigned(0 downto 0);
signal layer0_node48_MUX_bit_math_h_l546_c3_b0f6_iftrue : unsigned(7 downto 0);
signal layer0_node48_MUX_bit_math_h_l546_c3_b0f6_iffalse : unsigned(7 downto 0);
signal layer0_node48_MUX_bit_math_h_l546_c3_b0f6_return_output : unsigned(7 downto 0);

-- layer0_node49_MUX[bit_math_h_l557_c3_adcc]
signal layer0_node49_MUX_bit_math_h_l557_c3_adcc_cond : unsigned(0 downto 0);
signal layer0_node49_MUX_bit_math_h_l557_c3_adcc_iftrue : unsigned(7 downto 0);
signal layer0_node49_MUX_bit_math_h_l557_c3_adcc_iffalse : unsigned(7 downto 0);
signal layer0_node49_MUX_bit_math_h_l557_c3_adcc_return_output : unsigned(7 downto 0);

-- layer0_node50_MUX[bit_math_h_l568_c3_e90e]
signal layer0_node50_MUX_bit_math_h_l568_c3_e90e_cond : unsigned(0 downto 0);
signal layer0_node50_MUX_bit_math_h_l568_c3_e90e_iftrue : unsigned(7 downto 0);
signal layer0_node50_MUX_bit_math_h_l568_c3_e90e_iffalse : unsigned(7 downto 0);
signal layer0_node50_MUX_bit_math_h_l568_c3_e90e_return_output : unsigned(7 downto 0);

-- layer0_node51_MUX[bit_math_h_l579_c3_221f]
signal layer0_node51_MUX_bit_math_h_l579_c3_221f_cond : unsigned(0 downto 0);
signal layer0_node51_MUX_bit_math_h_l579_c3_221f_iftrue : unsigned(7 downto 0);
signal layer0_node51_MUX_bit_math_h_l579_c3_221f_iffalse : unsigned(7 downto 0);
signal layer0_node51_MUX_bit_math_h_l579_c3_221f_return_output : unsigned(7 downto 0);

-- layer0_node52_MUX[bit_math_h_l590_c3_70e0]
signal layer0_node52_MUX_bit_math_h_l590_c3_70e0_cond : unsigned(0 downto 0);
signal layer0_node52_MUX_bit_math_h_l590_c3_70e0_iftrue : unsigned(7 downto 0);
signal layer0_node52_MUX_bit_math_h_l590_c3_70e0_iffalse : unsigned(7 downto 0);
signal layer0_node52_MUX_bit_math_h_l590_c3_70e0_return_output : unsigned(7 downto 0);

-- layer0_node53_MUX[bit_math_h_l601_c3_e235]
signal layer0_node53_MUX_bit_math_h_l601_c3_e235_cond : unsigned(0 downto 0);
signal layer0_node53_MUX_bit_math_h_l601_c3_e235_iftrue : unsigned(7 downto 0);
signal layer0_node53_MUX_bit_math_h_l601_c3_e235_iffalse : unsigned(7 downto 0);
signal layer0_node53_MUX_bit_math_h_l601_c3_e235_return_output : unsigned(7 downto 0);

-- layer0_node54_MUX[bit_math_h_l612_c3_f982]
signal layer0_node54_MUX_bit_math_h_l612_c3_f982_cond : unsigned(0 downto 0);
signal layer0_node54_MUX_bit_math_h_l612_c3_f982_iftrue : unsigned(7 downto 0);
signal layer0_node54_MUX_bit_math_h_l612_c3_f982_iffalse : unsigned(7 downto 0);
signal layer0_node54_MUX_bit_math_h_l612_c3_f982_return_output : unsigned(7 downto 0);

-- layer0_node55_MUX[bit_math_h_l623_c3_bc3d]
signal layer0_node55_MUX_bit_math_h_l623_c3_bc3d_cond : unsigned(0 downto 0);
signal layer0_node55_MUX_bit_math_h_l623_c3_bc3d_iftrue : unsigned(7 downto 0);
signal layer0_node55_MUX_bit_math_h_l623_c3_bc3d_iffalse : unsigned(7 downto 0);
signal layer0_node55_MUX_bit_math_h_l623_c3_bc3d_return_output : unsigned(7 downto 0);

-- layer0_node56_MUX[bit_math_h_l634_c3_8e72]
signal layer0_node56_MUX_bit_math_h_l634_c3_8e72_cond : unsigned(0 downto 0);
signal layer0_node56_MUX_bit_math_h_l634_c3_8e72_iftrue : unsigned(7 downto 0);
signal layer0_node56_MUX_bit_math_h_l634_c3_8e72_iffalse : unsigned(7 downto 0);
signal layer0_node56_MUX_bit_math_h_l634_c3_8e72_return_output : unsigned(7 downto 0);

-- layer0_node57_MUX[bit_math_h_l645_c3_0789]
signal layer0_node57_MUX_bit_math_h_l645_c3_0789_cond : unsigned(0 downto 0);
signal layer0_node57_MUX_bit_math_h_l645_c3_0789_iftrue : unsigned(7 downto 0);
signal layer0_node57_MUX_bit_math_h_l645_c3_0789_iffalse : unsigned(7 downto 0);
signal layer0_node57_MUX_bit_math_h_l645_c3_0789_return_output : unsigned(7 downto 0);

-- layer0_node58_MUX[bit_math_h_l656_c3_d346]
signal layer0_node58_MUX_bit_math_h_l656_c3_d346_cond : unsigned(0 downto 0);
signal layer0_node58_MUX_bit_math_h_l656_c3_d346_iftrue : unsigned(7 downto 0);
signal layer0_node58_MUX_bit_math_h_l656_c3_d346_iffalse : unsigned(7 downto 0);
signal layer0_node58_MUX_bit_math_h_l656_c3_d346_return_output : unsigned(7 downto 0);

-- layer0_node59_MUX[bit_math_h_l667_c3_d31e]
signal layer0_node59_MUX_bit_math_h_l667_c3_d31e_cond : unsigned(0 downto 0);
signal layer0_node59_MUX_bit_math_h_l667_c3_d31e_iftrue : unsigned(7 downto 0);
signal layer0_node59_MUX_bit_math_h_l667_c3_d31e_iffalse : unsigned(7 downto 0);
signal layer0_node59_MUX_bit_math_h_l667_c3_d31e_return_output : unsigned(7 downto 0);

-- layer0_node60_MUX[bit_math_h_l678_c3_e120]
signal layer0_node60_MUX_bit_math_h_l678_c3_e120_cond : unsigned(0 downto 0);
signal layer0_node60_MUX_bit_math_h_l678_c3_e120_iftrue : unsigned(7 downto 0);
signal layer0_node60_MUX_bit_math_h_l678_c3_e120_iffalse : unsigned(7 downto 0);
signal layer0_node60_MUX_bit_math_h_l678_c3_e120_return_output : unsigned(7 downto 0);

-- layer0_node61_MUX[bit_math_h_l689_c3_a1a2]
signal layer0_node61_MUX_bit_math_h_l689_c3_a1a2_cond : unsigned(0 downto 0);
signal layer0_node61_MUX_bit_math_h_l689_c3_a1a2_iftrue : unsigned(7 downto 0);
signal layer0_node61_MUX_bit_math_h_l689_c3_a1a2_iffalse : unsigned(7 downto 0);
signal layer0_node61_MUX_bit_math_h_l689_c3_a1a2_return_output : unsigned(7 downto 0);

-- layer0_node62_MUX[bit_math_h_l700_c3_4595]
signal layer0_node62_MUX_bit_math_h_l700_c3_4595_cond : unsigned(0 downto 0);
signal layer0_node62_MUX_bit_math_h_l700_c3_4595_iftrue : unsigned(7 downto 0);
signal layer0_node62_MUX_bit_math_h_l700_c3_4595_iffalse : unsigned(7 downto 0);
signal layer0_node62_MUX_bit_math_h_l700_c3_4595_return_output : unsigned(7 downto 0);

-- layer0_node63_MUX[bit_math_h_l711_c3_c6ab]
signal layer0_node63_MUX_bit_math_h_l711_c3_c6ab_cond : unsigned(0 downto 0);
signal layer0_node63_MUX_bit_math_h_l711_c3_c6ab_iftrue : unsigned(7 downto 0);
signal layer0_node63_MUX_bit_math_h_l711_c3_c6ab_iffalse : unsigned(7 downto 0);
signal layer0_node63_MUX_bit_math_h_l711_c3_c6ab_return_output : unsigned(7 downto 0);

-- layer1_node0_MUX[bit_math_h_l728_c3_4268]
signal layer1_node0_MUX_bit_math_h_l728_c3_4268_cond : unsigned(0 downto 0);
signal layer1_node0_MUX_bit_math_h_l728_c3_4268_iftrue : unsigned(7 downto 0);
signal layer1_node0_MUX_bit_math_h_l728_c3_4268_iffalse : unsigned(7 downto 0);
signal layer1_node0_MUX_bit_math_h_l728_c3_4268_return_output : unsigned(7 downto 0);

-- layer1_node1_MUX[bit_math_h_l739_c3_ff28]
signal layer1_node1_MUX_bit_math_h_l739_c3_ff28_cond : unsigned(0 downto 0);
signal layer1_node1_MUX_bit_math_h_l739_c3_ff28_iftrue : unsigned(7 downto 0);
signal layer1_node1_MUX_bit_math_h_l739_c3_ff28_iffalse : unsigned(7 downto 0);
signal layer1_node1_MUX_bit_math_h_l739_c3_ff28_return_output : unsigned(7 downto 0);

-- layer1_node2_MUX[bit_math_h_l750_c3_543f]
signal layer1_node2_MUX_bit_math_h_l750_c3_543f_cond : unsigned(0 downto 0);
signal layer1_node2_MUX_bit_math_h_l750_c3_543f_iftrue : unsigned(7 downto 0);
signal layer1_node2_MUX_bit_math_h_l750_c3_543f_iffalse : unsigned(7 downto 0);
signal layer1_node2_MUX_bit_math_h_l750_c3_543f_return_output : unsigned(7 downto 0);

-- layer1_node3_MUX[bit_math_h_l761_c3_5c18]
signal layer1_node3_MUX_bit_math_h_l761_c3_5c18_cond : unsigned(0 downto 0);
signal layer1_node3_MUX_bit_math_h_l761_c3_5c18_iftrue : unsigned(7 downto 0);
signal layer1_node3_MUX_bit_math_h_l761_c3_5c18_iffalse : unsigned(7 downto 0);
signal layer1_node3_MUX_bit_math_h_l761_c3_5c18_return_output : unsigned(7 downto 0);

-- layer1_node4_MUX[bit_math_h_l772_c3_a66b]
signal layer1_node4_MUX_bit_math_h_l772_c3_a66b_cond : unsigned(0 downto 0);
signal layer1_node4_MUX_bit_math_h_l772_c3_a66b_iftrue : unsigned(7 downto 0);
signal layer1_node4_MUX_bit_math_h_l772_c3_a66b_iffalse : unsigned(7 downto 0);
signal layer1_node4_MUX_bit_math_h_l772_c3_a66b_return_output : unsigned(7 downto 0);

-- layer1_node5_MUX[bit_math_h_l783_c3_6db3]
signal layer1_node5_MUX_bit_math_h_l783_c3_6db3_cond : unsigned(0 downto 0);
signal layer1_node5_MUX_bit_math_h_l783_c3_6db3_iftrue : unsigned(7 downto 0);
signal layer1_node5_MUX_bit_math_h_l783_c3_6db3_iffalse : unsigned(7 downto 0);
signal layer1_node5_MUX_bit_math_h_l783_c3_6db3_return_output : unsigned(7 downto 0);

-- layer1_node6_MUX[bit_math_h_l794_c3_4c59]
signal layer1_node6_MUX_bit_math_h_l794_c3_4c59_cond : unsigned(0 downto 0);
signal layer1_node6_MUX_bit_math_h_l794_c3_4c59_iftrue : unsigned(7 downto 0);
signal layer1_node6_MUX_bit_math_h_l794_c3_4c59_iffalse : unsigned(7 downto 0);
signal layer1_node6_MUX_bit_math_h_l794_c3_4c59_return_output : unsigned(7 downto 0);

-- layer1_node7_MUX[bit_math_h_l805_c3_502f]
signal layer1_node7_MUX_bit_math_h_l805_c3_502f_cond : unsigned(0 downto 0);
signal layer1_node7_MUX_bit_math_h_l805_c3_502f_iftrue : unsigned(7 downto 0);
signal layer1_node7_MUX_bit_math_h_l805_c3_502f_iffalse : unsigned(7 downto 0);
signal layer1_node7_MUX_bit_math_h_l805_c3_502f_return_output : unsigned(7 downto 0);

-- layer1_node8_MUX[bit_math_h_l816_c3_1eec]
signal layer1_node8_MUX_bit_math_h_l816_c3_1eec_cond : unsigned(0 downto 0);
signal layer1_node8_MUX_bit_math_h_l816_c3_1eec_iftrue : unsigned(7 downto 0);
signal layer1_node8_MUX_bit_math_h_l816_c3_1eec_iffalse : unsigned(7 downto 0);
signal layer1_node8_MUX_bit_math_h_l816_c3_1eec_return_output : unsigned(7 downto 0);

-- layer1_node9_MUX[bit_math_h_l827_c3_d105]
signal layer1_node9_MUX_bit_math_h_l827_c3_d105_cond : unsigned(0 downto 0);
signal layer1_node9_MUX_bit_math_h_l827_c3_d105_iftrue : unsigned(7 downto 0);
signal layer1_node9_MUX_bit_math_h_l827_c3_d105_iffalse : unsigned(7 downto 0);
signal layer1_node9_MUX_bit_math_h_l827_c3_d105_return_output : unsigned(7 downto 0);

-- layer1_node10_MUX[bit_math_h_l838_c3_8a99]
signal layer1_node10_MUX_bit_math_h_l838_c3_8a99_cond : unsigned(0 downto 0);
signal layer1_node10_MUX_bit_math_h_l838_c3_8a99_iftrue : unsigned(7 downto 0);
signal layer1_node10_MUX_bit_math_h_l838_c3_8a99_iffalse : unsigned(7 downto 0);
signal layer1_node10_MUX_bit_math_h_l838_c3_8a99_return_output : unsigned(7 downto 0);

-- layer1_node11_MUX[bit_math_h_l849_c3_e0a5]
signal layer1_node11_MUX_bit_math_h_l849_c3_e0a5_cond : unsigned(0 downto 0);
signal layer1_node11_MUX_bit_math_h_l849_c3_e0a5_iftrue : unsigned(7 downto 0);
signal layer1_node11_MUX_bit_math_h_l849_c3_e0a5_iffalse : unsigned(7 downto 0);
signal layer1_node11_MUX_bit_math_h_l849_c3_e0a5_return_output : unsigned(7 downto 0);

-- layer1_node12_MUX[bit_math_h_l860_c3_53b9]
signal layer1_node12_MUX_bit_math_h_l860_c3_53b9_cond : unsigned(0 downto 0);
signal layer1_node12_MUX_bit_math_h_l860_c3_53b9_iftrue : unsigned(7 downto 0);
signal layer1_node12_MUX_bit_math_h_l860_c3_53b9_iffalse : unsigned(7 downto 0);
signal layer1_node12_MUX_bit_math_h_l860_c3_53b9_return_output : unsigned(7 downto 0);

-- layer1_node13_MUX[bit_math_h_l871_c3_672a]
signal layer1_node13_MUX_bit_math_h_l871_c3_672a_cond : unsigned(0 downto 0);
signal layer1_node13_MUX_bit_math_h_l871_c3_672a_iftrue : unsigned(7 downto 0);
signal layer1_node13_MUX_bit_math_h_l871_c3_672a_iffalse : unsigned(7 downto 0);
signal layer1_node13_MUX_bit_math_h_l871_c3_672a_return_output : unsigned(7 downto 0);

-- layer1_node14_MUX[bit_math_h_l882_c3_2725]
signal layer1_node14_MUX_bit_math_h_l882_c3_2725_cond : unsigned(0 downto 0);
signal layer1_node14_MUX_bit_math_h_l882_c3_2725_iftrue : unsigned(7 downto 0);
signal layer1_node14_MUX_bit_math_h_l882_c3_2725_iffalse : unsigned(7 downto 0);
signal layer1_node14_MUX_bit_math_h_l882_c3_2725_return_output : unsigned(7 downto 0);

-- layer1_node15_MUX[bit_math_h_l893_c3_b457]
signal layer1_node15_MUX_bit_math_h_l893_c3_b457_cond : unsigned(0 downto 0);
signal layer1_node15_MUX_bit_math_h_l893_c3_b457_iftrue : unsigned(7 downto 0);
signal layer1_node15_MUX_bit_math_h_l893_c3_b457_iffalse : unsigned(7 downto 0);
signal layer1_node15_MUX_bit_math_h_l893_c3_b457_return_output : unsigned(7 downto 0);

-- layer1_node16_MUX[bit_math_h_l904_c3_8832]
signal layer1_node16_MUX_bit_math_h_l904_c3_8832_cond : unsigned(0 downto 0);
signal layer1_node16_MUX_bit_math_h_l904_c3_8832_iftrue : unsigned(7 downto 0);
signal layer1_node16_MUX_bit_math_h_l904_c3_8832_iffalse : unsigned(7 downto 0);
signal layer1_node16_MUX_bit_math_h_l904_c3_8832_return_output : unsigned(7 downto 0);

-- layer1_node17_MUX[bit_math_h_l915_c3_0128]
signal layer1_node17_MUX_bit_math_h_l915_c3_0128_cond : unsigned(0 downto 0);
signal layer1_node17_MUX_bit_math_h_l915_c3_0128_iftrue : unsigned(7 downto 0);
signal layer1_node17_MUX_bit_math_h_l915_c3_0128_iffalse : unsigned(7 downto 0);
signal layer1_node17_MUX_bit_math_h_l915_c3_0128_return_output : unsigned(7 downto 0);

-- layer1_node18_MUX[bit_math_h_l926_c3_a8cf]
signal layer1_node18_MUX_bit_math_h_l926_c3_a8cf_cond : unsigned(0 downto 0);
signal layer1_node18_MUX_bit_math_h_l926_c3_a8cf_iftrue : unsigned(7 downto 0);
signal layer1_node18_MUX_bit_math_h_l926_c3_a8cf_iffalse : unsigned(7 downto 0);
signal layer1_node18_MUX_bit_math_h_l926_c3_a8cf_return_output : unsigned(7 downto 0);

-- layer1_node19_MUX[bit_math_h_l937_c3_3d6b]
signal layer1_node19_MUX_bit_math_h_l937_c3_3d6b_cond : unsigned(0 downto 0);
signal layer1_node19_MUX_bit_math_h_l937_c3_3d6b_iftrue : unsigned(7 downto 0);
signal layer1_node19_MUX_bit_math_h_l937_c3_3d6b_iffalse : unsigned(7 downto 0);
signal layer1_node19_MUX_bit_math_h_l937_c3_3d6b_return_output : unsigned(7 downto 0);

-- layer1_node20_MUX[bit_math_h_l948_c3_331f]
signal layer1_node20_MUX_bit_math_h_l948_c3_331f_cond : unsigned(0 downto 0);
signal layer1_node20_MUX_bit_math_h_l948_c3_331f_iftrue : unsigned(7 downto 0);
signal layer1_node20_MUX_bit_math_h_l948_c3_331f_iffalse : unsigned(7 downto 0);
signal layer1_node20_MUX_bit_math_h_l948_c3_331f_return_output : unsigned(7 downto 0);

-- layer1_node21_MUX[bit_math_h_l959_c3_32d5]
signal layer1_node21_MUX_bit_math_h_l959_c3_32d5_cond : unsigned(0 downto 0);
signal layer1_node21_MUX_bit_math_h_l959_c3_32d5_iftrue : unsigned(7 downto 0);
signal layer1_node21_MUX_bit_math_h_l959_c3_32d5_iffalse : unsigned(7 downto 0);
signal layer1_node21_MUX_bit_math_h_l959_c3_32d5_return_output : unsigned(7 downto 0);

-- layer1_node22_MUX[bit_math_h_l970_c3_56f9]
signal layer1_node22_MUX_bit_math_h_l970_c3_56f9_cond : unsigned(0 downto 0);
signal layer1_node22_MUX_bit_math_h_l970_c3_56f9_iftrue : unsigned(7 downto 0);
signal layer1_node22_MUX_bit_math_h_l970_c3_56f9_iffalse : unsigned(7 downto 0);
signal layer1_node22_MUX_bit_math_h_l970_c3_56f9_return_output : unsigned(7 downto 0);

-- layer1_node23_MUX[bit_math_h_l981_c3_251b]
signal layer1_node23_MUX_bit_math_h_l981_c3_251b_cond : unsigned(0 downto 0);
signal layer1_node23_MUX_bit_math_h_l981_c3_251b_iftrue : unsigned(7 downto 0);
signal layer1_node23_MUX_bit_math_h_l981_c3_251b_iffalse : unsigned(7 downto 0);
signal layer1_node23_MUX_bit_math_h_l981_c3_251b_return_output : unsigned(7 downto 0);

-- layer1_node24_MUX[bit_math_h_l992_c3_a508]
signal layer1_node24_MUX_bit_math_h_l992_c3_a508_cond : unsigned(0 downto 0);
signal layer1_node24_MUX_bit_math_h_l992_c3_a508_iftrue : unsigned(7 downto 0);
signal layer1_node24_MUX_bit_math_h_l992_c3_a508_iffalse : unsigned(7 downto 0);
signal layer1_node24_MUX_bit_math_h_l992_c3_a508_return_output : unsigned(7 downto 0);

-- layer1_node25_MUX[bit_math_h_l1003_c3_6bb3]
signal layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_cond : unsigned(0 downto 0);
signal layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_iftrue : unsigned(7 downto 0);
signal layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_iffalse : unsigned(7 downto 0);
signal layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_return_output : unsigned(7 downto 0);

-- layer1_node26_MUX[bit_math_h_l1014_c3_5bdb]
signal layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_cond : unsigned(0 downto 0);
signal layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_iftrue : unsigned(7 downto 0);
signal layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_iffalse : unsigned(7 downto 0);
signal layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_return_output : unsigned(7 downto 0);

-- layer1_node27_MUX[bit_math_h_l1025_c3_a0dc]
signal layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_cond : unsigned(0 downto 0);
signal layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_iftrue : unsigned(7 downto 0);
signal layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_iffalse : unsigned(7 downto 0);
signal layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_return_output : unsigned(7 downto 0);

-- layer1_node28_MUX[bit_math_h_l1036_c3_064f]
signal layer1_node28_MUX_bit_math_h_l1036_c3_064f_cond : unsigned(0 downto 0);
signal layer1_node28_MUX_bit_math_h_l1036_c3_064f_iftrue : unsigned(7 downto 0);
signal layer1_node28_MUX_bit_math_h_l1036_c3_064f_iffalse : unsigned(7 downto 0);
signal layer1_node28_MUX_bit_math_h_l1036_c3_064f_return_output : unsigned(7 downto 0);

-- layer1_node29_MUX[bit_math_h_l1047_c3_e950]
signal layer1_node29_MUX_bit_math_h_l1047_c3_e950_cond : unsigned(0 downto 0);
signal layer1_node29_MUX_bit_math_h_l1047_c3_e950_iftrue : unsigned(7 downto 0);
signal layer1_node29_MUX_bit_math_h_l1047_c3_e950_iffalse : unsigned(7 downto 0);
signal layer1_node29_MUX_bit_math_h_l1047_c3_e950_return_output : unsigned(7 downto 0);

-- layer1_node30_MUX[bit_math_h_l1058_c3_fdae]
signal layer1_node30_MUX_bit_math_h_l1058_c3_fdae_cond : unsigned(0 downto 0);
signal layer1_node30_MUX_bit_math_h_l1058_c3_fdae_iftrue : unsigned(7 downto 0);
signal layer1_node30_MUX_bit_math_h_l1058_c3_fdae_iffalse : unsigned(7 downto 0);
signal layer1_node30_MUX_bit_math_h_l1058_c3_fdae_return_output : unsigned(7 downto 0);

-- layer1_node31_MUX[bit_math_h_l1069_c3_6030]
signal layer1_node31_MUX_bit_math_h_l1069_c3_6030_cond : unsigned(0 downto 0);
signal layer1_node31_MUX_bit_math_h_l1069_c3_6030_iftrue : unsigned(7 downto 0);
signal layer1_node31_MUX_bit_math_h_l1069_c3_6030_iffalse : unsigned(7 downto 0);
signal layer1_node31_MUX_bit_math_h_l1069_c3_6030_return_output : unsigned(7 downto 0);

-- layer2_node0_MUX[bit_math_h_l1086_c3_122d]
signal layer2_node0_MUX_bit_math_h_l1086_c3_122d_cond : unsigned(0 downto 0);
signal layer2_node0_MUX_bit_math_h_l1086_c3_122d_iftrue : unsigned(7 downto 0);
signal layer2_node0_MUX_bit_math_h_l1086_c3_122d_iffalse : unsigned(7 downto 0);
signal layer2_node0_MUX_bit_math_h_l1086_c3_122d_return_output : unsigned(7 downto 0);

-- layer2_node1_MUX[bit_math_h_l1097_c3_fcc7]
signal layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_cond : unsigned(0 downto 0);
signal layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_iftrue : unsigned(7 downto 0);
signal layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_iffalse : unsigned(7 downto 0);
signal layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_return_output : unsigned(7 downto 0);

-- layer2_node2_MUX[bit_math_h_l1108_c3_b1b3]
signal layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_cond : unsigned(0 downto 0);
signal layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_iftrue : unsigned(7 downto 0);
signal layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_iffalse : unsigned(7 downto 0);
signal layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_return_output : unsigned(7 downto 0);

-- layer2_node3_MUX[bit_math_h_l1119_c3_946d]
signal layer2_node3_MUX_bit_math_h_l1119_c3_946d_cond : unsigned(0 downto 0);
signal layer2_node3_MUX_bit_math_h_l1119_c3_946d_iftrue : unsigned(7 downto 0);
signal layer2_node3_MUX_bit_math_h_l1119_c3_946d_iffalse : unsigned(7 downto 0);
signal layer2_node3_MUX_bit_math_h_l1119_c3_946d_return_output : unsigned(7 downto 0);

-- layer2_node4_MUX[bit_math_h_l1130_c3_1f93]
signal layer2_node4_MUX_bit_math_h_l1130_c3_1f93_cond : unsigned(0 downto 0);
signal layer2_node4_MUX_bit_math_h_l1130_c3_1f93_iftrue : unsigned(7 downto 0);
signal layer2_node4_MUX_bit_math_h_l1130_c3_1f93_iffalse : unsigned(7 downto 0);
signal layer2_node4_MUX_bit_math_h_l1130_c3_1f93_return_output : unsigned(7 downto 0);

-- layer2_node5_MUX[bit_math_h_l1141_c3_1425]
signal layer2_node5_MUX_bit_math_h_l1141_c3_1425_cond : unsigned(0 downto 0);
signal layer2_node5_MUX_bit_math_h_l1141_c3_1425_iftrue : unsigned(7 downto 0);
signal layer2_node5_MUX_bit_math_h_l1141_c3_1425_iffalse : unsigned(7 downto 0);
signal layer2_node5_MUX_bit_math_h_l1141_c3_1425_return_output : unsigned(7 downto 0);

-- layer2_node6_MUX[bit_math_h_l1152_c3_008a]
signal layer2_node6_MUX_bit_math_h_l1152_c3_008a_cond : unsigned(0 downto 0);
signal layer2_node6_MUX_bit_math_h_l1152_c3_008a_iftrue : unsigned(7 downto 0);
signal layer2_node6_MUX_bit_math_h_l1152_c3_008a_iffalse : unsigned(7 downto 0);
signal layer2_node6_MUX_bit_math_h_l1152_c3_008a_return_output : unsigned(7 downto 0);

-- layer2_node7_MUX[bit_math_h_l1163_c3_5ba0]
signal layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_cond : unsigned(0 downto 0);
signal layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_iftrue : unsigned(7 downto 0);
signal layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_iffalse : unsigned(7 downto 0);
signal layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_return_output : unsigned(7 downto 0);

-- layer2_node8_MUX[bit_math_h_l1174_c3_f1cf]
signal layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_cond : unsigned(0 downto 0);
signal layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_iftrue : unsigned(7 downto 0);
signal layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_iffalse : unsigned(7 downto 0);
signal layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_return_output : unsigned(7 downto 0);

-- layer2_node9_MUX[bit_math_h_l1185_c3_98c3]
signal layer2_node9_MUX_bit_math_h_l1185_c3_98c3_cond : unsigned(0 downto 0);
signal layer2_node9_MUX_bit_math_h_l1185_c3_98c3_iftrue : unsigned(7 downto 0);
signal layer2_node9_MUX_bit_math_h_l1185_c3_98c3_iffalse : unsigned(7 downto 0);
signal layer2_node9_MUX_bit_math_h_l1185_c3_98c3_return_output : unsigned(7 downto 0);

-- layer2_node10_MUX[bit_math_h_l1196_c3_1666]
signal layer2_node10_MUX_bit_math_h_l1196_c3_1666_cond : unsigned(0 downto 0);
signal layer2_node10_MUX_bit_math_h_l1196_c3_1666_iftrue : unsigned(7 downto 0);
signal layer2_node10_MUX_bit_math_h_l1196_c3_1666_iffalse : unsigned(7 downto 0);
signal layer2_node10_MUX_bit_math_h_l1196_c3_1666_return_output : unsigned(7 downto 0);

-- layer2_node11_MUX[bit_math_h_l1207_c3_b8de]
signal layer2_node11_MUX_bit_math_h_l1207_c3_b8de_cond : unsigned(0 downto 0);
signal layer2_node11_MUX_bit_math_h_l1207_c3_b8de_iftrue : unsigned(7 downto 0);
signal layer2_node11_MUX_bit_math_h_l1207_c3_b8de_iffalse : unsigned(7 downto 0);
signal layer2_node11_MUX_bit_math_h_l1207_c3_b8de_return_output : unsigned(7 downto 0);

-- layer2_node12_MUX[bit_math_h_l1218_c3_d8dc]
signal layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_cond : unsigned(0 downto 0);
signal layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_iftrue : unsigned(7 downto 0);
signal layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_iffalse : unsigned(7 downto 0);
signal layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_return_output : unsigned(7 downto 0);

-- layer2_node13_MUX[bit_math_h_l1229_c3_d585]
signal layer2_node13_MUX_bit_math_h_l1229_c3_d585_cond : unsigned(0 downto 0);
signal layer2_node13_MUX_bit_math_h_l1229_c3_d585_iftrue : unsigned(7 downto 0);
signal layer2_node13_MUX_bit_math_h_l1229_c3_d585_iffalse : unsigned(7 downto 0);
signal layer2_node13_MUX_bit_math_h_l1229_c3_d585_return_output : unsigned(7 downto 0);

-- layer2_node14_MUX[bit_math_h_l1240_c3_beb5]
signal layer2_node14_MUX_bit_math_h_l1240_c3_beb5_cond : unsigned(0 downto 0);
signal layer2_node14_MUX_bit_math_h_l1240_c3_beb5_iftrue : unsigned(7 downto 0);
signal layer2_node14_MUX_bit_math_h_l1240_c3_beb5_iffalse : unsigned(7 downto 0);
signal layer2_node14_MUX_bit_math_h_l1240_c3_beb5_return_output : unsigned(7 downto 0);

-- layer2_node15_MUX[bit_math_h_l1251_c3_7550]
signal layer2_node15_MUX_bit_math_h_l1251_c3_7550_cond : unsigned(0 downto 0);
signal layer2_node15_MUX_bit_math_h_l1251_c3_7550_iftrue : unsigned(7 downto 0);
signal layer2_node15_MUX_bit_math_h_l1251_c3_7550_iffalse : unsigned(7 downto 0);
signal layer2_node15_MUX_bit_math_h_l1251_c3_7550_return_output : unsigned(7 downto 0);

-- layer3_node0_MUX[bit_math_h_l1268_c3_302d]
signal layer3_node0_MUX_bit_math_h_l1268_c3_302d_cond : unsigned(0 downto 0);
signal layer3_node0_MUX_bit_math_h_l1268_c3_302d_iftrue : unsigned(7 downto 0);
signal layer3_node0_MUX_bit_math_h_l1268_c3_302d_iffalse : unsigned(7 downto 0);
signal layer3_node0_MUX_bit_math_h_l1268_c3_302d_return_output : unsigned(7 downto 0);

-- layer3_node1_MUX[bit_math_h_l1279_c3_fd3b]
signal layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_cond : unsigned(0 downto 0);
signal layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_iftrue : unsigned(7 downto 0);
signal layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_iffalse : unsigned(7 downto 0);
signal layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_return_output : unsigned(7 downto 0);

-- layer3_node2_MUX[bit_math_h_l1290_c3_5e3f]
signal layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_cond : unsigned(0 downto 0);
signal layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_iftrue : unsigned(7 downto 0);
signal layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_iffalse : unsigned(7 downto 0);
signal layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_return_output : unsigned(7 downto 0);

-- layer3_node3_MUX[bit_math_h_l1301_c3_84c3]
signal layer3_node3_MUX_bit_math_h_l1301_c3_84c3_cond : unsigned(0 downto 0);
signal layer3_node3_MUX_bit_math_h_l1301_c3_84c3_iftrue : unsigned(7 downto 0);
signal layer3_node3_MUX_bit_math_h_l1301_c3_84c3_iffalse : unsigned(7 downto 0);
signal layer3_node3_MUX_bit_math_h_l1301_c3_84c3_return_output : unsigned(7 downto 0);

-- layer3_node4_MUX[bit_math_h_l1312_c3_8c96]
signal layer3_node4_MUX_bit_math_h_l1312_c3_8c96_cond : unsigned(0 downto 0);
signal layer3_node4_MUX_bit_math_h_l1312_c3_8c96_iftrue : unsigned(7 downto 0);
signal layer3_node4_MUX_bit_math_h_l1312_c3_8c96_iffalse : unsigned(7 downto 0);
signal layer3_node4_MUX_bit_math_h_l1312_c3_8c96_return_output : unsigned(7 downto 0);

-- layer3_node5_MUX[bit_math_h_l1323_c3_57ee]
signal layer3_node5_MUX_bit_math_h_l1323_c3_57ee_cond : unsigned(0 downto 0);
signal layer3_node5_MUX_bit_math_h_l1323_c3_57ee_iftrue : unsigned(7 downto 0);
signal layer3_node5_MUX_bit_math_h_l1323_c3_57ee_iffalse : unsigned(7 downto 0);
signal layer3_node5_MUX_bit_math_h_l1323_c3_57ee_return_output : unsigned(7 downto 0);

-- layer3_node6_MUX[bit_math_h_l1334_c3_f24c]
signal layer3_node6_MUX_bit_math_h_l1334_c3_f24c_cond : unsigned(0 downto 0);
signal layer3_node6_MUX_bit_math_h_l1334_c3_f24c_iftrue : unsigned(7 downto 0);
signal layer3_node6_MUX_bit_math_h_l1334_c3_f24c_iffalse : unsigned(7 downto 0);
signal layer3_node6_MUX_bit_math_h_l1334_c3_f24c_return_output : unsigned(7 downto 0);

-- layer3_node7_MUX[bit_math_h_l1345_c3_c68c]
signal layer3_node7_MUX_bit_math_h_l1345_c3_c68c_cond : unsigned(0 downto 0);
signal layer3_node7_MUX_bit_math_h_l1345_c3_c68c_iftrue : unsigned(7 downto 0);
signal layer3_node7_MUX_bit_math_h_l1345_c3_c68c_iffalse : unsigned(7 downto 0);
signal layer3_node7_MUX_bit_math_h_l1345_c3_c68c_return_output : unsigned(7 downto 0);

-- layer4_node0_MUX[bit_math_h_l1362_c3_a122]
signal layer4_node0_MUX_bit_math_h_l1362_c3_a122_cond : unsigned(0 downto 0);
signal layer4_node0_MUX_bit_math_h_l1362_c3_a122_iftrue : unsigned(7 downto 0);
signal layer4_node0_MUX_bit_math_h_l1362_c3_a122_iffalse : unsigned(7 downto 0);
signal layer4_node0_MUX_bit_math_h_l1362_c3_a122_return_output : unsigned(7 downto 0);

-- layer4_node1_MUX[bit_math_h_l1373_c3_c86f]
signal layer4_node1_MUX_bit_math_h_l1373_c3_c86f_cond : unsigned(0 downto 0);
signal layer4_node1_MUX_bit_math_h_l1373_c3_c86f_iftrue : unsigned(7 downto 0);
signal layer4_node1_MUX_bit_math_h_l1373_c3_c86f_iffalse : unsigned(7 downto 0);
signal layer4_node1_MUX_bit_math_h_l1373_c3_c86f_return_output : unsigned(7 downto 0);

-- layer4_node2_MUX[bit_math_h_l1384_c3_76f0]
signal layer4_node2_MUX_bit_math_h_l1384_c3_76f0_cond : unsigned(0 downto 0);
signal layer4_node2_MUX_bit_math_h_l1384_c3_76f0_iftrue : unsigned(7 downto 0);
signal layer4_node2_MUX_bit_math_h_l1384_c3_76f0_iffalse : unsigned(7 downto 0);
signal layer4_node2_MUX_bit_math_h_l1384_c3_76f0_return_output : unsigned(7 downto 0);

-- layer4_node3_MUX[bit_math_h_l1395_c3_5649]
signal layer4_node3_MUX_bit_math_h_l1395_c3_5649_cond : unsigned(0 downto 0);
signal layer4_node3_MUX_bit_math_h_l1395_c3_5649_iftrue : unsigned(7 downto 0);
signal layer4_node3_MUX_bit_math_h_l1395_c3_5649_iffalse : unsigned(7 downto 0);
signal layer4_node3_MUX_bit_math_h_l1395_c3_5649_return_output : unsigned(7 downto 0);

-- layer5_node0_MUX[bit_math_h_l1412_c3_c6a2]
signal layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_cond : unsigned(0 downto 0);
signal layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_iftrue : unsigned(7 downto 0);
signal layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_iffalse : unsigned(7 downto 0);
signal layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_return_output : unsigned(7 downto 0);

-- layer5_node1_MUX[bit_math_h_l1423_c3_d92a]
signal layer5_node1_MUX_bit_math_h_l1423_c3_d92a_cond : unsigned(0 downto 0);
signal layer5_node1_MUX_bit_math_h_l1423_c3_d92a_iftrue : unsigned(7 downto 0);
signal layer5_node1_MUX_bit_math_h_l1423_c3_d92a_iffalse : unsigned(7 downto 0);
signal layer5_node1_MUX_bit_math_h_l1423_c3_d92a_return_output : unsigned(7 downto 0);

-- layer6_node0_MUX[bit_math_h_l1440_c3_43c9]
signal layer6_node0_MUX_bit_math_h_l1440_c3_43c9_cond : unsigned(0 downto 0);
signal layer6_node0_MUX_bit_math_h_l1440_c3_43c9_iftrue : unsigned(7 downto 0);
signal layer6_node0_MUX_bit_math_h_l1440_c3_43c9_iffalse : unsigned(7 downto 0);
signal layer6_node0_MUX_bit_math_h_l1440_c3_43c9_return_output : unsigned(7 downto 0);

function uint7_0_0( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(0- i);
      end loop;
return return_output;
end function;

function uint7_1_1( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(1- i);
      end loop;
return return_output;
end function;

function uint7_2_2( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(2- i);
      end loop;
return return_output;
end function;

function uint7_3_3( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(3- i);
      end loop;
return return_output;
end function;

function uint7_4_4( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(4- i);
      end loop;
return return_output;
end function;

function uint7_5_5( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(5- i);
      end loop;
return return_output;
end function;

function uint7_6_6( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(6- i);
      end loop;
return return_output;
end function;


begin

-- SUBMODULE INSTANCES 
-- layer0_node0_MUX_bit_math_h_l18_c3_ce9b
layer0_node0_MUX_bit_math_h_l18_c3_ce9b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node0_MUX_bit_math_h_l18_c3_ce9b_cond,
layer0_node0_MUX_bit_math_h_l18_c3_ce9b_iftrue,
layer0_node0_MUX_bit_math_h_l18_c3_ce9b_iffalse,
layer0_node0_MUX_bit_math_h_l18_c3_ce9b_return_output);

-- layer0_node1_MUX_bit_math_h_l29_c3_0e94
layer0_node1_MUX_bit_math_h_l29_c3_0e94 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node1_MUX_bit_math_h_l29_c3_0e94_cond,
layer0_node1_MUX_bit_math_h_l29_c3_0e94_iftrue,
layer0_node1_MUX_bit_math_h_l29_c3_0e94_iffalse,
layer0_node1_MUX_bit_math_h_l29_c3_0e94_return_output);

-- layer0_node2_MUX_bit_math_h_l40_c3_e2d9
layer0_node2_MUX_bit_math_h_l40_c3_e2d9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node2_MUX_bit_math_h_l40_c3_e2d9_cond,
layer0_node2_MUX_bit_math_h_l40_c3_e2d9_iftrue,
layer0_node2_MUX_bit_math_h_l40_c3_e2d9_iffalse,
layer0_node2_MUX_bit_math_h_l40_c3_e2d9_return_output);

-- layer0_node3_MUX_bit_math_h_l51_c3_edc9
layer0_node3_MUX_bit_math_h_l51_c3_edc9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node3_MUX_bit_math_h_l51_c3_edc9_cond,
layer0_node3_MUX_bit_math_h_l51_c3_edc9_iftrue,
layer0_node3_MUX_bit_math_h_l51_c3_edc9_iffalse,
layer0_node3_MUX_bit_math_h_l51_c3_edc9_return_output);

-- layer0_node4_MUX_bit_math_h_l62_c3_f389
layer0_node4_MUX_bit_math_h_l62_c3_f389 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node4_MUX_bit_math_h_l62_c3_f389_cond,
layer0_node4_MUX_bit_math_h_l62_c3_f389_iftrue,
layer0_node4_MUX_bit_math_h_l62_c3_f389_iffalse,
layer0_node4_MUX_bit_math_h_l62_c3_f389_return_output);

-- layer0_node5_MUX_bit_math_h_l73_c3_d655
layer0_node5_MUX_bit_math_h_l73_c3_d655 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node5_MUX_bit_math_h_l73_c3_d655_cond,
layer0_node5_MUX_bit_math_h_l73_c3_d655_iftrue,
layer0_node5_MUX_bit_math_h_l73_c3_d655_iffalse,
layer0_node5_MUX_bit_math_h_l73_c3_d655_return_output);

-- layer0_node6_MUX_bit_math_h_l84_c3_5cd3
layer0_node6_MUX_bit_math_h_l84_c3_5cd3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node6_MUX_bit_math_h_l84_c3_5cd3_cond,
layer0_node6_MUX_bit_math_h_l84_c3_5cd3_iftrue,
layer0_node6_MUX_bit_math_h_l84_c3_5cd3_iffalse,
layer0_node6_MUX_bit_math_h_l84_c3_5cd3_return_output);

-- layer0_node7_MUX_bit_math_h_l95_c3_5030
layer0_node7_MUX_bit_math_h_l95_c3_5030 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node7_MUX_bit_math_h_l95_c3_5030_cond,
layer0_node7_MUX_bit_math_h_l95_c3_5030_iftrue,
layer0_node7_MUX_bit_math_h_l95_c3_5030_iffalse,
layer0_node7_MUX_bit_math_h_l95_c3_5030_return_output);

-- layer0_node8_MUX_bit_math_h_l106_c3_32cb
layer0_node8_MUX_bit_math_h_l106_c3_32cb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node8_MUX_bit_math_h_l106_c3_32cb_cond,
layer0_node8_MUX_bit_math_h_l106_c3_32cb_iftrue,
layer0_node8_MUX_bit_math_h_l106_c3_32cb_iffalse,
layer0_node8_MUX_bit_math_h_l106_c3_32cb_return_output);

-- layer0_node9_MUX_bit_math_h_l117_c3_4b42
layer0_node9_MUX_bit_math_h_l117_c3_4b42 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node9_MUX_bit_math_h_l117_c3_4b42_cond,
layer0_node9_MUX_bit_math_h_l117_c3_4b42_iftrue,
layer0_node9_MUX_bit_math_h_l117_c3_4b42_iffalse,
layer0_node9_MUX_bit_math_h_l117_c3_4b42_return_output);

-- layer0_node10_MUX_bit_math_h_l128_c3_06f3
layer0_node10_MUX_bit_math_h_l128_c3_06f3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node10_MUX_bit_math_h_l128_c3_06f3_cond,
layer0_node10_MUX_bit_math_h_l128_c3_06f3_iftrue,
layer0_node10_MUX_bit_math_h_l128_c3_06f3_iffalse,
layer0_node10_MUX_bit_math_h_l128_c3_06f3_return_output);

-- layer0_node11_MUX_bit_math_h_l139_c3_dbfc
layer0_node11_MUX_bit_math_h_l139_c3_dbfc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node11_MUX_bit_math_h_l139_c3_dbfc_cond,
layer0_node11_MUX_bit_math_h_l139_c3_dbfc_iftrue,
layer0_node11_MUX_bit_math_h_l139_c3_dbfc_iffalse,
layer0_node11_MUX_bit_math_h_l139_c3_dbfc_return_output);

-- layer0_node12_MUX_bit_math_h_l150_c3_6613
layer0_node12_MUX_bit_math_h_l150_c3_6613 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node12_MUX_bit_math_h_l150_c3_6613_cond,
layer0_node12_MUX_bit_math_h_l150_c3_6613_iftrue,
layer0_node12_MUX_bit_math_h_l150_c3_6613_iffalse,
layer0_node12_MUX_bit_math_h_l150_c3_6613_return_output);

-- layer0_node13_MUX_bit_math_h_l161_c3_fd42
layer0_node13_MUX_bit_math_h_l161_c3_fd42 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node13_MUX_bit_math_h_l161_c3_fd42_cond,
layer0_node13_MUX_bit_math_h_l161_c3_fd42_iftrue,
layer0_node13_MUX_bit_math_h_l161_c3_fd42_iffalse,
layer0_node13_MUX_bit_math_h_l161_c3_fd42_return_output);

-- layer0_node14_MUX_bit_math_h_l172_c3_154a
layer0_node14_MUX_bit_math_h_l172_c3_154a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node14_MUX_bit_math_h_l172_c3_154a_cond,
layer0_node14_MUX_bit_math_h_l172_c3_154a_iftrue,
layer0_node14_MUX_bit_math_h_l172_c3_154a_iffalse,
layer0_node14_MUX_bit_math_h_l172_c3_154a_return_output);

-- layer0_node15_MUX_bit_math_h_l183_c3_5274
layer0_node15_MUX_bit_math_h_l183_c3_5274 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node15_MUX_bit_math_h_l183_c3_5274_cond,
layer0_node15_MUX_bit_math_h_l183_c3_5274_iftrue,
layer0_node15_MUX_bit_math_h_l183_c3_5274_iffalse,
layer0_node15_MUX_bit_math_h_l183_c3_5274_return_output);

-- layer0_node16_MUX_bit_math_h_l194_c3_7a7d
layer0_node16_MUX_bit_math_h_l194_c3_7a7d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node16_MUX_bit_math_h_l194_c3_7a7d_cond,
layer0_node16_MUX_bit_math_h_l194_c3_7a7d_iftrue,
layer0_node16_MUX_bit_math_h_l194_c3_7a7d_iffalse,
layer0_node16_MUX_bit_math_h_l194_c3_7a7d_return_output);

-- layer0_node17_MUX_bit_math_h_l205_c3_42ac
layer0_node17_MUX_bit_math_h_l205_c3_42ac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node17_MUX_bit_math_h_l205_c3_42ac_cond,
layer0_node17_MUX_bit_math_h_l205_c3_42ac_iftrue,
layer0_node17_MUX_bit_math_h_l205_c3_42ac_iffalse,
layer0_node17_MUX_bit_math_h_l205_c3_42ac_return_output);

-- layer0_node18_MUX_bit_math_h_l216_c3_b8f1
layer0_node18_MUX_bit_math_h_l216_c3_b8f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node18_MUX_bit_math_h_l216_c3_b8f1_cond,
layer0_node18_MUX_bit_math_h_l216_c3_b8f1_iftrue,
layer0_node18_MUX_bit_math_h_l216_c3_b8f1_iffalse,
layer0_node18_MUX_bit_math_h_l216_c3_b8f1_return_output);

-- layer0_node19_MUX_bit_math_h_l227_c3_0b12
layer0_node19_MUX_bit_math_h_l227_c3_0b12 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node19_MUX_bit_math_h_l227_c3_0b12_cond,
layer0_node19_MUX_bit_math_h_l227_c3_0b12_iftrue,
layer0_node19_MUX_bit_math_h_l227_c3_0b12_iffalse,
layer0_node19_MUX_bit_math_h_l227_c3_0b12_return_output);

-- layer0_node20_MUX_bit_math_h_l238_c3_091e
layer0_node20_MUX_bit_math_h_l238_c3_091e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node20_MUX_bit_math_h_l238_c3_091e_cond,
layer0_node20_MUX_bit_math_h_l238_c3_091e_iftrue,
layer0_node20_MUX_bit_math_h_l238_c3_091e_iffalse,
layer0_node20_MUX_bit_math_h_l238_c3_091e_return_output);

-- layer0_node21_MUX_bit_math_h_l249_c3_44d2
layer0_node21_MUX_bit_math_h_l249_c3_44d2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node21_MUX_bit_math_h_l249_c3_44d2_cond,
layer0_node21_MUX_bit_math_h_l249_c3_44d2_iftrue,
layer0_node21_MUX_bit_math_h_l249_c3_44d2_iffalse,
layer0_node21_MUX_bit_math_h_l249_c3_44d2_return_output);

-- layer0_node22_MUX_bit_math_h_l260_c3_db28
layer0_node22_MUX_bit_math_h_l260_c3_db28 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node22_MUX_bit_math_h_l260_c3_db28_cond,
layer0_node22_MUX_bit_math_h_l260_c3_db28_iftrue,
layer0_node22_MUX_bit_math_h_l260_c3_db28_iffalse,
layer0_node22_MUX_bit_math_h_l260_c3_db28_return_output);

-- layer0_node23_MUX_bit_math_h_l271_c3_0038
layer0_node23_MUX_bit_math_h_l271_c3_0038 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node23_MUX_bit_math_h_l271_c3_0038_cond,
layer0_node23_MUX_bit_math_h_l271_c3_0038_iftrue,
layer0_node23_MUX_bit_math_h_l271_c3_0038_iffalse,
layer0_node23_MUX_bit_math_h_l271_c3_0038_return_output);

-- layer0_node24_MUX_bit_math_h_l282_c3_1d56
layer0_node24_MUX_bit_math_h_l282_c3_1d56 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node24_MUX_bit_math_h_l282_c3_1d56_cond,
layer0_node24_MUX_bit_math_h_l282_c3_1d56_iftrue,
layer0_node24_MUX_bit_math_h_l282_c3_1d56_iffalse,
layer0_node24_MUX_bit_math_h_l282_c3_1d56_return_output);

-- layer0_node25_MUX_bit_math_h_l293_c3_fa3c
layer0_node25_MUX_bit_math_h_l293_c3_fa3c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node25_MUX_bit_math_h_l293_c3_fa3c_cond,
layer0_node25_MUX_bit_math_h_l293_c3_fa3c_iftrue,
layer0_node25_MUX_bit_math_h_l293_c3_fa3c_iffalse,
layer0_node25_MUX_bit_math_h_l293_c3_fa3c_return_output);

-- layer0_node26_MUX_bit_math_h_l304_c3_220e
layer0_node26_MUX_bit_math_h_l304_c3_220e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node26_MUX_bit_math_h_l304_c3_220e_cond,
layer0_node26_MUX_bit_math_h_l304_c3_220e_iftrue,
layer0_node26_MUX_bit_math_h_l304_c3_220e_iffalse,
layer0_node26_MUX_bit_math_h_l304_c3_220e_return_output);

-- layer0_node27_MUX_bit_math_h_l315_c3_37d2
layer0_node27_MUX_bit_math_h_l315_c3_37d2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node27_MUX_bit_math_h_l315_c3_37d2_cond,
layer0_node27_MUX_bit_math_h_l315_c3_37d2_iftrue,
layer0_node27_MUX_bit_math_h_l315_c3_37d2_iffalse,
layer0_node27_MUX_bit_math_h_l315_c3_37d2_return_output);

-- layer0_node28_MUX_bit_math_h_l326_c3_af14
layer0_node28_MUX_bit_math_h_l326_c3_af14 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node28_MUX_bit_math_h_l326_c3_af14_cond,
layer0_node28_MUX_bit_math_h_l326_c3_af14_iftrue,
layer0_node28_MUX_bit_math_h_l326_c3_af14_iffalse,
layer0_node28_MUX_bit_math_h_l326_c3_af14_return_output);

-- layer0_node29_MUX_bit_math_h_l337_c3_d491
layer0_node29_MUX_bit_math_h_l337_c3_d491 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node29_MUX_bit_math_h_l337_c3_d491_cond,
layer0_node29_MUX_bit_math_h_l337_c3_d491_iftrue,
layer0_node29_MUX_bit_math_h_l337_c3_d491_iffalse,
layer0_node29_MUX_bit_math_h_l337_c3_d491_return_output);

-- layer0_node30_MUX_bit_math_h_l348_c3_46cf
layer0_node30_MUX_bit_math_h_l348_c3_46cf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node30_MUX_bit_math_h_l348_c3_46cf_cond,
layer0_node30_MUX_bit_math_h_l348_c3_46cf_iftrue,
layer0_node30_MUX_bit_math_h_l348_c3_46cf_iffalse,
layer0_node30_MUX_bit_math_h_l348_c3_46cf_return_output);

-- layer0_node31_MUX_bit_math_h_l359_c3_1ee6
layer0_node31_MUX_bit_math_h_l359_c3_1ee6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node31_MUX_bit_math_h_l359_c3_1ee6_cond,
layer0_node31_MUX_bit_math_h_l359_c3_1ee6_iftrue,
layer0_node31_MUX_bit_math_h_l359_c3_1ee6_iffalse,
layer0_node31_MUX_bit_math_h_l359_c3_1ee6_return_output);

-- layer0_node32_MUX_bit_math_h_l370_c3_ee39
layer0_node32_MUX_bit_math_h_l370_c3_ee39 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node32_MUX_bit_math_h_l370_c3_ee39_cond,
layer0_node32_MUX_bit_math_h_l370_c3_ee39_iftrue,
layer0_node32_MUX_bit_math_h_l370_c3_ee39_iffalse,
layer0_node32_MUX_bit_math_h_l370_c3_ee39_return_output);

-- layer0_node33_MUX_bit_math_h_l381_c3_f57d
layer0_node33_MUX_bit_math_h_l381_c3_f57d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node33_MUX_bit_math_h_l381_c3_f57d_cond,
layer0_node33_MUX_bit_math_h_l381_c3_f57d_iftrue,
layer0_node33_MUX_bit_math_h_l381_c3_f57d_iffalse,
layer0_node33_MUX_bit_math_h_l381_c3_f57d_return_output);

-- layer0_node34_MUX_bit_math_h_l392_c3_8d4e
layer0_node34_MUX_bit_math_h_l392_c3_8d4e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node34_MUX_bit_math_h_l392_c3_8d4e_cond,
layer0_node34_MUX_bit_math_h_l392_c3_8d4e_iftrue,
layer0_node34_MUX_bit_math_h_l392_c3_8d4e_iffalse,
layer0_node34_MUX_bit_math_h_l392_c3_8d4e_return_output);

-- layer0_node35_MUX_bit_math_h_l403_c3_fa1f
layer0_node35_MUX_bit_math_h_l403_c3_fa1f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node35_MUX_bit_math_h_l403_c3_fa1f_cond,
layer0_node35_MUX_bit_math_h_l403_c3_fa1f_iftrue,
layer0_node35_MUX_bit_math_h_l403_c3_fa1f_iffalse,
layer0_node35_MUX_bit_math_h_l403_c3_fa1f_return_output);

-- layer0_node36_MUX_bit_math_h_l414_c3_39b4
layer0_node36_MUX_bit_math_h_l414_c3_39b4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node36_MUX_bit_math_h_l414_c3_39b4_cond,
layer0_node36_MUX_bit_math_h_l414_c3_39b4_iftrue,
layer0_node36_MUX_bit_math_h_l414_c3_39b4_iffalse,
layer0_node36_MUX_bit_math_h_l414_c3_39b4_return_output);

-- layer0_node37_MUX_bit_math_h_l425_c3_3900
layer0_node37_MUX_bit_math_h_l425_c3_3900 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node37_MUX_bit_math_h_l425_c3_3900_cond,
layer0_node37_MUX_bit_math_h_l425_c3_3900_iftrue,
layer0_node37_MUX_bit_math_h_l425_c3_3900_iffalse,
layer0_node37_MUX_bit_math_h_l425_c3_3900_return_output);

-- layer0_node38_MUX_bit_math_h_l436_c3_bea2
layer0_node38_MUX_bit_math_h_l436_c3_bea2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node38_MUX_bit_math_h_l436_c3_bea2_cond,
layer0_node38_MUX_bit_math_h_l436_c3_bea2_iftrue,
layer0_node38_MUX_bit_math_h_l436_c3_bea2_iffalse,
layer0_node38_MUX_bit_math_h_l436_c3_bea2_return_output);

-- layer0_node39_MUX_bit_math_h_l447_c3_3acc
layer0_node39_MUX_bit_math_h_l447_c3_3acc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node39_MUX_bit_math_h_l447_c3_3acc_cond,
layer0_node39_MUX_bit_math_h_l447_c3_3acc_iftrue,
layer0_node39_MUX_bit_math_h_l447_c3_3acc_iffalse,
layer0_node39_MUX_bit_math_h_l447_c3_3acc_return_output);

-- layer0_node40_MUX_bit_math_h_l458_c3_f867
layer0_node40_MUX_bit_math_h_l458_c3_f867 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node40_MUX_bit_math_h_l458_c3_f867_cond,
layer0_node40_MUX_bit_math_h_l458_c3_f867_iftrue,
layer0_node40_MUX_bit_math_h_l458_c3_f867_iffalse,
layer0_node40_MUX_bit_math_h_l458_c3_f867_return_output);

-- layer0_node41_MUX_bit_math_h_l469_c3_2ffe
layer0_node41_MUX_bit_math_h_l469_c3_2ffe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node41_MUX_bit_math_h_l469_c3_2ffe_cond,
layer0_node41_MUX_bit_math_h_l469_c3_2ffe_iftrue,
layer0_node41_MUX_bit_math_h_l469_c3_2ffe_iffalse,
layer0_node41_MUX_bit_math_h_l469_c3_2ffe_return_output);

-- layer0_node42_MUX_bit_math_h_l480_c3_1c62
layer0_node42_MUX_bit_math_h_l480_c3_1c62 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node42_MUX_bit_math_h_l480_c3_1c62_cond,
layer0_node42_MUX_bit_math_h_l480_c3_1c62_iftrue,
layer0_node42_MUX_bit_math_h_l480_c3_1c62_iffalse,
layer0_node42_MUX_bit_math_h_l480_c3_1c62_return_output);

-- layer0_node43_MUX_bit_math_h_l491_c3_7943
layer0_node43_MUX_bit_math_h_l491_c3_7943 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node43_MUX_bit_math_h_l491_c3_7943_cond,
layer0_node43_MUX_bit_math_h_l491_c3_7943_iftrue,
layer0_node43_MUX_bit_math_h_l491_c3_7943_iffalse,
layer0_node43_MUX_bit_math_h_l491_c3_7943_return_output);

-- layer0_node44_MUX_bit_math_h_l502_c3_15dc
layer0_node44_MUX_bit_math_h_l502_c3_15dc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node44_MUX_bit_math_h_l502_c3_15dc_cond,
layer0_node44_MUX_bit_math_h_l502_c3_15dc_iftrue,
layer0_node44_MUX_bit_math_h_l502_c3_15dc_iffalse,
layer0_node44_MUX_bit_math_h_l502_c3_15dc_return_output);

-- layer0_node45_MUX_bit_math_h_l513_c3_d638
layer0_node45_MUX_bit_math_h_l513_c3_d638 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node45_MUX_bit_math_h_l513_c3_d638_cond,
layer0_node45_MUX_bit_math_h_l513_c3_d638_iftrue,
layer0_node45_MUX_bit_math_h_l513_c3_d638_iffalse,
layer0_node45_MUX_bit_math_h_l513_c3_d638_return_output);

-- layer0_node46_MUX_bit_math_h_l524_c3_fdc0
layer0_node46_MUX_bit_math_h_l524_c3_fdc0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node46_MUX_bit_math_h_l524_c3_fdc0_cond,
layer0_node46_MUX_bit_math_h_l524_c3_fdc0_iftrue,
layer0_node46_MUX_bit_math_h_l524_c3_fdc0_iffalse,
layer0_node46_MUX_bit_math_h_l524_c3_fdc0_return_output);

-- layer0_node47_MUX_bit_math_h_l535_c3_1640
layer0_node47_MUX_bit_math_h_l535_c3_1640 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node47_MUX_bit_math_h_l535_c3_1640_cond,
layer0_node47_MUX_bit_math_h_l535_c3_1640_iftrue,
layer0_node47_MUX_bit_math_h_l535_c3_1640_iffalse,
layer0_node47_MUX_bit_math_h_l535_c3_1640_return_output);

-- layer0_node48_MUX_bit_math_h_l546_c3_b0f6
layer0_node48_MUX_bit_math_h_l546_c3_b0f6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node48_MUX_bit_math_h_l546_c3_b0f6_cond,
layer0_node48_MUX_bit_math_h_l546_c3_b0f6_iftrue,
layer0_node48_MUX_bit_math_h_l546_c3_b0f6_iffalse,
layer0_node48_MUX_bit_math_h_l546_c3_b0f6_return_output);

-- layer0_node49_MUX_bit_math_h_l557_c3_adcc
layer0_node49_MUX_bit_math_h_l557_c3_adcc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node49_MUX_bit_math_h_l557_c3_adcc_cond,
layer0_node49_MUX_bit_math_h_l557_c3_adcc_iftrue,
layer0_node49_MUX_bit_math_h_l557_c3_adcc_iffalse,
layer0_node49_MUX_bit_math_h_l557_c3_adcc_return_output);

-- layer0_node50_MUX_bit_math_h_l568_c3_e90e
layer0_node50_MUX_bit_math_h_l568_c3_e90e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node50_MUX_bit_math_h_l568_c3_e90e_cond,
layer0_node50_MUX_bit_math_h_l568_c3_e90e_iftrue,
layer0_node50_MUX_bit_math_h_l568_c3_e90e_iffalse,
layer0_node50_MUX_bit_math_h_l568_c3_e90e_return_output);

-- layer0_node51_MUX_bit_math_h_l579_c3_221f
layer0_node51_MUX_bit_math_h_l579_c3_221f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node51_MUX_bit_math_h_l579_c3_221f_cond,
layer0_node51_MUX_bit_math_h_l579_c3_221f_iftrue,
layer0_node51_MUX_bit_math_h_l579_c3_221f_iffalse,
layer0_node51_MUX_bit_math_h_l579_c3_221f_return_output);

-- layer0_node52_MUX_bit_math_h_l590_c3_70e0
layer0_node52_MUX_bit_math_h_l590_c3_70e0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node52_MUX_bit_math_h_l590_c3_70e0_cond,
layer0_node52_MUX_bit_math_h_l590_c3_70e0_iftrue,
layer0_node52_MUX_bit_math_h_l590_c3_70e0_iffalse,
layer0_node52_MUX_bit_math_h_l590_c3_70e0_return_output);

-- layer0_node53_MUX_bit_math_h_l601_c3_e235
layer0_node53_MUX_bit_math_h_l601_c3_e235 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node53_MUX_bit_math_h_l601_c3_e235_cond,
layer0_node53_MUX_bit_math_h_l601_c3_e235_iftrue,
layer0_node53_MUX_bit_math_h_l601_c3_e235_iffalse,
layer0_node53_MUX_bit_math_h_l601_c3_e235_return_output);

-- layer0_node54_MUX_bit_math_h_l612_c3_f982
layer0_node54_MUX_bit_math_h_l612_c3_f982 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node54_MUX_bit_math_h_l612_c3_f982_cond,
layer0_node54_MUX_bit_math_h_l612_c3_f982_iftrue,
layer0_node54_MUX_bit_math_h_l612_c3_f982_iffalse,
layer0_node54_MUX_bit_math_h_l612_c3_f982_return_output);

-- layer0_node55_MUX_bit_math_h_l623_c3_bc3d
layer0_node55_MUX_bit_math_h_l623_c3_bc3d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node55_MUX_bit_math_h_l623_c3_bc3d_cond,
layer0_node55_MUX_bit_math_h_l623_c3_bc3d_iftrue,
layer0_node55_MUX_bit_math_h_l623_c3_bc3d_iffalse,
layer0_node55_MUX_bit_math_h_l623_c3_bc3d_return_output);

-- layer0_node56_MUX_bit_math_h_l634_c3_8e72
layer0_node56_MUX_bit_math_h_l634_c3_8e72 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node56_MUX_bit_math_h_l634_c3_8e72_cond,
layer0_node56_MUX_bit_math_h_l634_c3_8e72_iftrue,
layer0_node56_MUX_bit_math_h_l634_c3_8e72_iffalse,
layer0_node56_MUX_bit_math_h_l634_c3_8e72_return_output);

-- layer0_node57_MUX_bit_math_h_l645_c3_0789
layer0_node57_MUX_bit_math_h_l645_c3_0789 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node57_MUX_bit_math_h_l645_c3_0789_cond,
layer0_node57_MUX_bit_math_h_l645_c3_0789_iftrue,
layer0_node57_MUX_bit_math_h_l645_c3_0789_iffalse,
layer0_node57_MUX_bit_math_h_l645_c3_0789_return_output);

-- layer0_node58_MUX_bit_math_h_l656_c3_d346
layer0_node58_MUX_bit_math_h_l656_c3_d346 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node58_MUX_bit_math_h_l656_c3_d346_cond,
layer0_node58_MUX_bit_math_h_l656_c3_d346_iftrue,
layer0_node58_MUX_bit_math_h_l656_c3_d346_iffalse,
layer0_node58_MUX_bit_math_h_l656_c3_d346_return_output);

-- layer0_node59_MUX_bit_math_h_l667_c3_d31e
layer0_node59_MUX_bit_math_h_l667_c3_d31e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node59_MUX_bit_math_h_l667_c3_d31e_cond,
layer0_node59_MUX_bit_math_h_l667_c3_d31e_iftrue,
layer0_node59_MUX_bit_math_h_l667_c3_d31e_iffalse,
layer0_node59_MUX_bit_math_h_l667_c3_d31e_return_output);

-- layer0_node60_MUX_bit_math_h_l678_c3_e120
layer0_node60_MUX_bit_math_h_l678_c3_e120 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node60_MUX_bit_math_h_l678_c3_e120_cond,
layer0_node60_MUX_bit_math_h_l678_c3_e120_iftrue,
layer0_node60_MUX_bit_math_h_l678_c3_e120_iffalse,
layer0_node60_MUX_bit_math_h_l678_c3_e120_return_output);

-- layer0_node61_MUX_bit_math_h_l689_c3_a1a2
layer0_node61_MUX_bit_math_h_l689_c3_a1a2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node61_MUX_bit_math_h_l689_c3_a1a2_cond,
layer0_node61_MUX_bit_math_h_l689_c3_a1a2_iftrue,
layer0_node61_MUX_bit_math_h_l689_c3_a1a2_iffalse,
layer0_node61_MUX_bit_math_h_l689_c3_a1a2_return_output);

-- layer0_node62_MUX_bit_math_h_l700_c3_4595
layer0_node62_MUX_bit_math_h_l700_c3_4595 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node62_MUX_bit_math_h_l700_c3_4595_cond,
layer0_node62_MUX_bit_math_h_l700_c3_4595_iftrue,
layer0_node62_MUX_bit_math_h_l700_c3_4595_iffalse,
layer0_node62_MUX_bit_math_h_l700_c3_4595_return_output);

-- layer0_node63_MUX_bit_math_h_l711_c3_c6ab
layer0_node63_MUX_bit_math_h_l711_c3_c6ab : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node63_MUX_bit_math_h_l711_c3_c6ab_cond,
layer0_node63_MUX_bit_math_h_l711_c3_c6ab_iftrue,
layer0_node63_MUX_bit_math_h_l711_c3_c6ab_iffalse,
layer0_node63_MUX_bit_math_h_l711_c3_c6ab_return_output);

-- layer1_node0_MUX_bit_math_h_l728_c3_4268
layer1_node0_MUX_bit_math_h_l728_c3_4268 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node0_MUX_bit_math_h_l728_c3_4268_cond,
layer1_node0_MUX_bit_math_h_l728_c3_4268_iftrue,
layer1_node0_MUX_bit_math_h_l728_c3_4268_iffalse,
layer1_node0_MUX_bit_math_h_l728_c3_4268_return_output);

-- layer1_node1_MUX_bit_math_h_l739_c3_ff28
layer1_node1_MUX_bit_math_h_l739_c3_ff28 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node1_MUX_bit_math_h_l739_c3_ff28_cond,
layer1_node1_MUX_bit_math_h_l739_c3_ff28_iftrue,
layer1_node1_MUX_bit_math_h_l739_c3_ff28_iffalse,
layer1_node1_MUX_bit_math_h_l739_c3_ff28_return_output);

-- layer1_node2_MUX_bit_math_h_l750_c3_543f
layer1_node2_MUX_bit_math_h_l750_c3_543f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node2_MUX_bit_math_h_l750_c3_543f_cond,
layer1_node2_MUX_bit_math_h_l750_c3_543f_iftrue,
layer1_node2_MUX_bit_math_h_l750_c3_543f_iffalse,
layer1_node2_MUX_bit_math_h_l750_c3_543f_return_output);

-- layer1_node3_MUX_bit_math_h_l761_c3_5c18
layer1_node3_MUX_bit_math_h_l761_c3_5c18 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node3_MUX_bit_math_h_l761_c3_5c18_cond,
layer1_node3_MUX_bit_math_h_l761_c3_5c18_iftrue,
layer1_node3_MUX_bit_math_h_l761_c3_5c18_iffalse,
layer1_node3_MUX_bit_math_h_l761_c3_5c18_return_output);

-- layer1_node4_MUX_bit_math_h_l772_c3_a66b
layer1_node4_MUX_bit_math_h_l772_c3_a66b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node4_MUX_bit_math_h_l772_c3_a66b_cond,
layer1_node4_MUX_bit_math_h_l772_c3_a66b_iftrue,
layer1_node4_MUX_bit_math_h_l772_c3_a66b_iffalse,
layer1_node4_MUX_bit_math_h_l772_c3_a66b_return_output);

-- layer1_node5_MUX_bit_math_h_l783_c3_6db3
layer1_node5_MUX_bit_math_h_l783_c3_6db3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node5_MUX_bit_math_h_l783_c3_6db3_cond,
layer1_node5_MUX_bit_math_h_l783_c3_6db3_iftrue,
layer1_node5_MUX_bit_math_h_l783_c3_6db3_iffalse,
layer1_node5_MUX_bit_math_h_l783_c3_6db3_return_output);

-- layer1_node6_MUX_bit_math_h_l794_c3_4c59
layer1_node6_MUX_bit_math_h_l794_c3_4c59 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node6_MUX_bit_math_h_l794_c3_4c59_cond,
layer1_node6_MUX_bit_math_h_l794_c3_4c59_iftrue,
layer1_node6_MUX_bit_math_h_l794_c3_4c59_iffalse,
layer1_node6_MUX_bit_math_h_l794_c3_4c59_return_output);

-- layer1_node7_MUX_bit_math_h_l805_c3_502f
layer1_node7_MUX_bit_math_h_l805_c3_502f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node7_MUX_bit_math_h_l805_c3_502f_cond,
layer1_node7_MUX_bit_math_h_l805_c3_502f_iftrue,
layer1_node7_MUX_bit_math_h_l805_c3_502f_iffalse,
layer1_node7_MUX_bit_math_h_l805_c3_502f_return_output);

-- layer1_node8_MUX_bit_math_h_l816_c3_1eec
layer1_node8_MUX_bit_math_h_l816_c3_1eec : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node8_MUX_bit_math_h_l816_c3_1eec_cond,
layer1_node8_MUX_bit_math_h_l816_c3_1eec_iftrue,
layer1_node8_MUX_bit_math_h_l816_c3_1eec_iffalse,
layer1_node8_MUX_bit_math_h_l816_c3_1eec_return_output);

-- layer1_node9_MUX_bit_math_h_l827_c3_d105
layer1_node9_MUX_bit_math_h_l827_c3_d105 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node9_MUX_bit_math_h_l827_c3_d105_cond,
layer1_node9_MUX_bit_math_h_l827_c3_d105_iftrue,
layer1_node9_MUX_bit_math_h_l827_c3_d105_iffalse,
layer1_node9_MUX_bit_math_h_l827_c3_d105_return_output);

-- layer1_node10_MUX_bit_math_h_l838_c3_8a99
layer1_node10_MUX_bit_math_h_l838_c3_8a99 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node10_MUX_bit_math_h_l838_c3_8a99_cond,
layer1_node10_MUX_bit_math_h_l838_c3_8a99_iftrue,
layer1_node10_MUX_bit_math_h_l838_c3_8a99_iffalse,
layer1_node10_MUX_bit_math_h_l838_c3_8a99_return_output);

-- layer1_node11_MUX_bit_math_h_l849_c3_e0a5
layer1_node11_MUX_bit_math_h_l849_c3_e0a5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node11_MUX_bit_math_h_l849_c3_e0a5_cond,
layer1_node11_MUX_bit_math_h_l849_c3_e0a5_iftrue,
layer1_node11_MUX_bit_math_h_l849_c3_e0a5_iffalse,
layer1_node11_MUX_bit_math_h_l849_c3_e0a5_return_output);

-- layer1_node12_MUX_bit_math_h_l860_c3_53b9
layer1_node12_MUX_bit_math_h_l860_c3_53b9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node12_MUX_bit_math_h_l860_c3_53b9_cond,
layer1_node12_MUX_bit_math_h_l860_c3_53b9_iftrue,
layer1_node12_MUX_bit_math_h_l860_c3_53b9_iffalse,
layer1_node12_MUX_bit_math_h_l860_c3_53b9_return_output);

-- layer1_node13_MUX_bit_math_h_l871_c3_672a
layer1_node13_MUX_bit_math_h_l871_c3_672a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node13_MUX_bit_math_h_l871_c3_672a_cond,
layer1_node13_MUX_bit_math_h_l871_c3_672a_iftrue,
layer1_node13_MUX_bit_math_h_l871_c3_672a_iffalse,
layer1_node13_MUX_bit_math_h_l871_c3_672a_return_output);

-- layer1_node14_MUX_bit_math_h_l882_c3_2725
layer1_node14_MUX_bit_math_h_l882_c3_2725 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node14_MUX_bit_math_h_l882_c3_2725_cond,
layer1_node14_MUX_bit_math_h_l882_c3_2725_iftrue,
layer1_node14_MUX_bit_math_h_l882_c3_2725_iffalse,
layer1_node14_MUX_bit_math_h_l882_c3_2725_return_output);

-- layer1_node15_MUX_bit_math_h_l893_c3_b457
layer1_node15_MUX_bit_math_h_l893_c3_b457 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node15_MUX_bit_math_h_l893_c3_b457_cond,
layer1_node15_MUX_bit_math_h_l893_c3_b457_iftrue,
layer1_node15_MUX_bit_math_h_l893_c3_b457_iffalse,
layer1_node15_MUX_bit_math_h_l893_c3_b457_return_output);

-- layer1_node16_MUX_bit_math_h_l904_c3_8832
layer1_node16_MUX_bit_math_h_l904_c3_8832 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node16_MUX_bit_math_h_l904_c3_8832_cond,
layer1_node16_MUX_bit_math_h_l904_c3_8832_iftrue,
layer1_node16_MUX_bit_math_h_l904_c3_8832_iffalse,
layer1_node16_MUX_bit_math_h_l904_c3_8832_return_output);

-- layer1_node17_MUX_bit_math_h_l915_c3_0128
layer1_node17_MUX_bit_math_h_l915_c3_0128 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node17_MUX_bit_math_h_l915_c3_0128_cond,
layer1_node17_MUX_bit_math_h_l915_c3_0128_iftrue,
layer1_node17_MUX_bit_math_h_l915_c3_0128_iffalse,
layer1_node17_MUX_bit_math_h_l915_c3_0128_return_output);

-- layer1_node18_MUX_bit_math_h_l926_c3_a8cf
layer1_node18_MUX_bit_math_h_l926_c3_a8cf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node18_MUX_bit_math_h_l926_c3_a8cf_cond,
layer1_node18_MUX_bit_math_h_l926_c3_a8cf_iftrue,
layer1_node18_MUX_bit_math_h_l926_c3_a8cf_iffalse,
layer1_node18_MUX_bit_math_h_l926_c3_a8cf_return_output);

-- layer1_node19_MUX_bit_math_h_l937_c3_3d6b
layer1_node19_MUX_bit_math_h_l937_c3_3d6b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node19_MUX_bit_math_h_l937_c3_3d6b_cond,
layer1_node19_MUX_bit_math_h_l937_c3_3d6b_iftrue,
layer1_node19_MUX_bit_math_h_l937_c3_3d6b_iffalse,
layer1_node19_MUX_bit_math_h_l937_c3_3d6b_return_output);

-- layer1_node20_MUX_bit_math_h_l948_c3_331f
layer1_node20_MUX_bit_math_h_l948_c3_331f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node20_MUX_bit_math_h_l948_c3_331f_cond,
layer1_node20_MUX_bit_math_h_l948_c3_331f_iftrue,
layer1_node20_MUX_bit_math_h_l948_c3_331f_iffalse,
layer1_node20_MUX_bit_math_h_l948_c3_331f_return_output);

-- layer1_node21_MUX_bit_math_h_l959_c3_32d5
layer1_node21_MUX_bit_math_h_l959_c3_32d5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node21_MUX_bit_math_h_l959_c3_32d5_cond,
layer1_node21_MUX_bit_math_h_l959_c3_32d5_iftrue,
layer1_node21_MUX_bit_math_h_l959_c3_32d5_iffalse,
layer1_node21_MUX_bit_math_h_l959_c3_32d5_return_output);

-- layer1_node22_MUX_bit_math_h_l970_c3_56f9
layer1_node22_MUX_bit_math_h_l970_c3_56f9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node22_MUX_bit_math_h_l970_c3_56f9_cond,
layer1_node22_MUX_bit_math_h_l970_c3_56f9_iftrue,
layer1_node22_MUX_bit_math_h_l970_c3_56f9_iffalse,
layer1_node22_MUX_bit_math_h_l970_c3_56f9_return_output);

-- layer1_node23_MUX_bit_math_h_l981_c3_251b
layer1_node23_MUX_bit_math_h_l981_c3_251b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node23_MUX_bit_math_h_l981_c3_251b_cond,
layer1_node23_MUX_bit_math_h_l981_c3_251b_iftrue,
layer1_node23_MUX_bit_math_h_l981_c3_251b_iffalse,
layer1_node23_MUX_bit_math_h_l981_c3_251b_return_output);

-- layer1_node24_MUX_bit_math_h_l992_c3_a508
layer1_node24_MUX_bit_math_h_l992_c3_a508 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node24_MUX_bit_math_h_l992_c3_a508_cond,
layer1_node24_MUX_bit_math_h_l992_c3_a508_iftrue,
layer1_node24_MUX_bit_math_h_l992_c3_a508_iffalse,
layer1_node24_MUX_bit_math_h_l992_c3_a508_return_output);

-- layer1_node25_MUX_bit_math_h_l1003_c3_6bb3
layer1_node25_MUX_bit_math_h_l1003_c3_6bb3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_cond,
layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_iftrue,
layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_iffalse,
layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_return_output);

-- layer1_node26_MUX_bit_math_h_l1014_c3_5bdb
layer1_node26_MUX_bit_math_h_l1014_c3_5bdb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_cond,
layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_iftrue,
layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_iffalse,
layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_return_output);

-- layer1_node27_MUX_bit_math_h_l1025_c3_a0dc
layer1_node27_MUX_bit_math_h_l1025_c3_a0dc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_cond,
layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_iftrue,
layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_iffalse,
layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_return_output);

-- layer1_node28_MUX_bit_math_h_l1036_c3_064f
layer1_node28_MUX_bit_math_h_l1036_c3_064f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node28_MUX_bit_math_h_l1036_c3_064f_cond,
layer1_node28_MUX_bit_math_h_l1036_c3_064f_iftrue,
layer1_node28_MUX_bit_math_h_l1036_c3_064f_iffalse,
layer1_node28_MUX_bit_math_h_l1036_c3_064f_return_output);

-- layer1_node29_MUX_bit_math_h_l1047_c3_e950
layer1_node29_MUX_bit_math_h_l1047_c3_e950 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node29_MUX_bit_math_h_l1047_c3_e950_cond,
layer1_node29_MUX_bit_math_h_l1047_c3_e950_iftrue,
layer1_node29_MUX_bit_math_h_l1047_c3_e950_iffalse,
layer1_node29_MUX_bit_math_h_l1047_c3_e950_return_output);

-- layer1_node30_MUX_bit_math_h_l1058_c3_fdae
layer1_node30_MUX_bit_math_h_l1058_c3_fdae : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node30_MUX_bit_math_h_l1058_c3_fdae_cond,
layer1_node30_MUX_bit_math_h_l1058_c3_fdae_iftrue,
layer1_node30_MUX_bit_math_h_l1058_c3_fdae_iffalse,
layer1_node30_MUX_bit_math_h_l1058_c3_fdae_return_output);

-- layer1_node31_MUX_bit_math_h_l1069_c3_6030
layer1_node31_MUX_bit_math_h_l1069_c3_6030 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node31_MUX_bit_math_h_l1069_c3_6030_cond,
layer1_node31_MUX_bit_math_h_l1069_c3_6030_iftrue,
layer1_node31_MUX_bit_math_h_l1069_c3_6030_iffalse,
layer1_node31_MUX_bit_math_h_l1069_c3_6030_return_output);

-- layer2_node0_MUX_bit_math_h_l1086_c3_122d
layer2_node0_MUX_bit_math_h_l1086_c3_122d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node0_MUX_bit_math_h_l1086_c3_122d_cond,
layer2_node0_MUX_bit_math_h_l1086_c3_122d_iftrue,
layer2_node0_MUX_bit_math_h_l1086_c3_122d_iffalse,
layer2_node0_MUX_bit_math_h_l1086_c3_122d_return_output);

-- layer2_node1_MUX_bit_math_h_l1097_c3_fcc7
layer2_node1_MUX_bit_math_h_l1097_c3_fcc7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_cond,
layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_iftrue,
layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_iffalse,
layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_return_output);

-- layer2_node2_MUX_bit_math_h_l1108_c3_b1b3
layer2_node2_MUX_bit_math_h_l1108_c3_b1b3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_cond,
layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_iftrue,
layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_iffalse,
layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_return_output);

-- layer2_node3_MUX_bit_math_h_l1119_c3_946d
layer2_node3_MUX_bit_math_h_l1119_c3_946d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node3_MUX_bit_math_h_l1119_c3_946d_cond,
layer2_node3_MUX_bit_math_h_l1119_c3_946d_iftrue,
layer2_node3_MUX_bit_math_h_l1119_c3_946d_iffalse,
layer2_node3_MUX_bit_math_h_l1119_c3_946d_return_output);

-- layer2_node4_MUX_bit_math_h_l1130_c3_1f93
layer2_node4_MUX_bit_math_h_l1130_c3_1f93 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node4_MUX_bit_math_h_l1130_c3_1f93_cond,
layer2_node4_MUX_bit_math_h_l1130_c3_1f93_iftrue,
layer2_node4_MUX_bit_math_h_l1130_c3_1f93_iffalse,
layer2_node4_MUX_bit_math_h_l1130_c3_1f93_return_output);

-- layer2_node5_MUX_bit_math_h_l1141_c3_1425
layer2_node5_MUX_bit_math_h_l1141_c3_1425 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node5_MUX_bit_math_h_l1141_c3_1425_cond,
layer2_node5_MUX_bit_math_h_l1141_c3_1425_iftrue,
layer2_node5_MUX_bit_math_h_l1141_c3_1425_iffalse,
layer2_node5_MUX_bit_math_h_l1141_c3_1425_return_output);

-- layer2_node6_MUX_bit_math_h_l1152_c3_008a
layer2_node6_MUX_bit_math_h_l1152_c3_008a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node6_MUX_bit_math_h_l1152_c3_008a_cond,
layer2_node6_MUX_bit_math_h_l1152_c3_008a_iftrue,
layer2_node6_MUX_bit_math_h_l1152_c3_008a_iffalse,
layer2_node6_MUX_bit_math_h_l1152_c3_008a_return_output);

-- layer2_node7_MUX_bit_math_h_l1163_c3_5ba0
layer2_node7_MUX_bit_math_h_l1163_c3_5ba0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_cond,
layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_iftrue,
layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_iffalse,
layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_return_output);

-- layer2_node8_MUX_bit_math_h_l1174_c3_f1cf
layer2_node8_MUX_bit_math_h_l1174_c3_f1cf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_cond,
layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_iftrue,
layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_iffalse,
layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_return_output);

-- layer2_node9_MUX_bit_math_h_l1185_c3_98c3
layer2_node9_MUX_bit_math_h_l1185_c3_98c3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node9_MUX_bit_math_h_l1185_c3_98c3_cond,
layer2_node9_MUX_bit_math_h_l1185_c3_98c3_iftrue,
layer2_node9_MUX_bit_math_h_l1185_c3_98c3_iffalse,
layer2_node9_MUX_bit_math_h_l1185_c3_98c3_return_output);

-- layer2_node10_MUX_bit_math_h_l1196_c3_1666
layer2_node10_MUX_bit_math_h_l1196_c3_1666 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node10_MUX_bit_math_h_l1196_c3_1666_cond,
layer2_node10_MUX_bit_math_h_l1196_c3_1666_iftrue,
layer2_node10_MUX_bit_math_h_l1196_c3_1666_iffalse,
layer2_node10_MUX_bit_math_h_l1196_c3_1666_return_output);

-- layer2_node11_MUX_bit_math_h_l1207_c3_b8de
layer2_node11_MUX_bit_math_h_l1207_c3_b8de : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node11_MUX_bit_math_h_l1207_c3_b8de_cond,
layer2_node11_MUX_bit_math_h_l1207_c3_b8de_iftrue,
layer2_node11_MUX_bit_math_h_l1207_c3_b8de_iffalse,
layer2_node11_MUX_bit_math_h_l1207_c3_b8de_return_output);

-- layer2_node12_MUX_bit_math_h_l1218_c3_d8dc
layer2_node12_MUX_bit_math_h_l1218_c3_d8dc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_cond,
layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_iftrue,
layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_iffalse,
layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_return_output);

-- layer2_node13_MUX_bit_math_h_l1229_c3_d585
layer2_node13_MUX_bit_math_h_l1229_c3_d585 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node13_MUX_bit_math_h_l1229_c3_d585_cond,
layer2_node13_MUX_bit_math_h_l1229_c3_d585_iftrue,
layer2_node13_MUX_bit_math_h_l1229_c3_d585_iffalse,
layer2_node13_MUX_bit_math_h_l1229_c3_d585_return_output);

-- layer2_node14_MUX_bit_math_h_l1240_c3_beb5
layer2_node14_MUX_bit_math_h_l1240_c3_beb5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node14_MUX_bit_math_h_l1240_c3_beb5_cond,
layer2_node14_MUX_bit_math_h_l1240_c3_beb5_iftrue,
layer2_node14_MUX_bit_math_h_l1240_c3_beb5_iffalse,
layer2_node14_MUX_bit_math_h_l1240_c3_beb5_return_output);

-- layer2_node15_MUX_bit_math_h_l1251_c3_7550
layer2_node15_MUX_bit_math_h_l1251_c3_7550 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node15_MUX_bit_math_h_l1251_c3_7550_cond,
layer2_node15_MUX_bit_math_h_l1251_c3_7550_iftrue,
layer2_node15_MUX_bit_math_h_l1251_c3_7550_iffalse,
layer2_node15_MUX_bit_math_h_l1251_c3_7550_return_output);

-- layer3_node0_MUX_bit_math_h_l1268_c3_302d
layer3_node0_MUX_bit_math_h_l1268_c3_302d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node0_MUX_bit_math_h_l1268_c3_302d_cond,
layer3_node0_MUX_bit_math_h_l1268_c3_302d_iftrue,
layer3_node0_MUX_bit_math_h_l1268_c3_302d_iffalse,
layer3_node0_MUX_bit_math_h_l1268_c3_302d_return_output);

-- layer3_node1_MUX_bit_math_h_l1279_c3_fd3b
layer3_node1_MUX_bit_math_h_l1279_c3_fd3b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_cond,
layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_iftrue,
layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_iffalse,
layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_return_output);

-- layer3_node2_MUX_bit_math_h_l1290_c3_5e3f
layer3_node2_MUX_bit_math_h_l1290_c3_5e3f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_cond,
layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_iftrue,
layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_iffalse,
layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_return_output);

-- layer3_node3_MUX_bit_math_h_l1301_c3_84c3
layer3_node3_MUX_bit_math_h_l1301_c3_84c3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node3_MUX_bit_math_h_l1301_c3_84c3_cond,
layer3_node3_MUX_bit_math_h_l1301_c3_84c3_iftrue,
layer3_node3_MUX_bit_math_h_l1301_c3_84c3_iffalse,
layer3_node3_MUX_bit_math_h_l1301_c3_84c3_return_output);

-- layer3_node4_MUX_bit_math_h_l1312_c3_8c96
layer3_node4_MUX_bit_math_h_l1312_c3_8c96 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node4_MUX_bit_math_h_l1312_c3_8c96_cond,
layer3_node4_MUX_bit_math_h_l1312_c3_8c96_iftrue,
layer3_node4_MUX_bit_math_h_l1312_c3_8c96_iffalse,
layer3_node4_MUX_bit_math_h_l1312_c3_8c96_return_output);

-- layer3_node5_MUX_bit_math_h_l1323_c3_57ee
layer3_node5_MUX_bit_math_h_l1323_c3_57ee : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node5_MUX_bit_math_h_l1323_c3_57ee_cond,
layer3_node5_MUX_bit_math_h_l1323_c3_57ee_iftrue,
layer3_node5_MUX_bit_math_h_l1323_c3_57ee_iffalse,
layer3_node5_MUX_bit_math_h_l1323_c3_57ee_return_output);

-- layer3_node6_MUX_bit_math_h_l1334_c3_f24c
layer3_node6_MUX_bit_math_h_l1334_c3_f24c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node6_MUX_bit_math_h_l1334_c3_f24c_cond,
layer3_node6_MUX_bit_math_h_l1334_c3_f24c_iftrue,
layer3_node6_MUX_bit_math_h_l1334_c3_f24c_iffalse,
layer3_node6_MUX_bit_math_h_l1334_c3_f24c_return_output);

-- layer3_node7_MUX_bit_math_h_l1345_c3_c68c
layer3_node7_MUX_bit_math_h_l1345_c3_c68c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node7_MUX_bit_math_h_l1345_c3_c68c_cond,
layer3_node7_MUX_bit_math_h_l1345_c3_c68c_iftrue,
layer3_node7_MUX_bit_math_h_l1345_c3_c68c_iffalse,
layer3_node7_MUX_bit_math_h_l1345_c3_c68c_return_output);

-- layer4_node0_MUX_bit_math_h_l1362_c3_a122
layer4_node0_MUX_bit_math_h_l1362_c3_a122 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer4_node0_MUX_bit_math_h_l1362_c3_a122_cond,
layer4_node0_MUX_bit_math_h_l1362_c3_a122_iftrue,
layer4_node0_MUX_bit_math_h_l1362_c3_a122_iffalse,
layer4_node0_MUX_bit_math_h_l1362_c3_a122_return_output);

-- layer4_node1_MUX_bit_math_h_l1373_c3_c86f
layer4_node1_MUX_bit_math_h_l1373_c3_c86f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer4_node1_MUX_bit_math_h_l1373_c3_c86f_cond,
layer4_node1_MUX_bit_math_h_l1373_c3_c86f_iftrue,
layer4_node1_MUX_bit_math_h_l1373_c3_c86f_iffalse,
layer4_node1_MUX_bit_math_h_l1373_c3_c86f_return_output);

-- layer4_node2_MUX_bit_math_h_l1384_c3_76f0
layer4_node2_MUX_bit_math_h_l1384_c3_76f0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer4_node2_MUX_bit_math_h_l1384_c3_76f0_cond,
layer4_node2_MUX_bit_math_h_l1384_c3_76f0_iftrue,
layer4_node2_MUX_bit_math_h_l1384_c3_76f0_iffalse,
layer4_node2_MUX_bit_math_h_l1384_c3_76f0_return_output);

-- layer4_node3_MUX_bit_math_h_l1395_c3_5649
layer4_node3_MUX_bit_math_h_l1395_c3_5649 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer4_node3_MUX_bit_math_h_l1395_c3_5649_cond,
layer4_node3_MUX_bit_math_h_l1395_c3_5649_iftrue,
layer4_node3_MUX_bit_math_h_l1395_c3_5649_iffalse,
layer4_node3_MUX_bit_math_h_l1395_c3_5649_return_output);

-- layer5_node0_MUX_bit_math_h_l1412_c3_c6a2
layer5_node0_MUX_bit_math_h_l1412_c3_c6a2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_cond,
layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_iftrue,
layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_iffalse,
layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_return_output);

-- layer5_node1_MUX_bit_math_h_l1423_c3_d92a
layer5_node1_MUX_bit_math_h_l1423_c3_d92a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer5_node1_MUX_bit_math_h_l1423_c3_d92a_cond,
layer5_node1_MUX_bit_math_h_l1423_c3_d92a_iftrue,
layer5_node1_MUX_bit_math_h_l1423_c3_d92a_iffalse,
layer5_node1_MUX_bit_math_h_l1423_c3_d92a_return_output);

-- layer6_node0_MUX_bit_math_h_l1440_c3_43c9
layer6_node0_MUX_bit_math_h_l1440_c3_43c9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer6_node0_MUX_bit_math_h_l1440_c3_43c9_cond,
layer6_node0_MUX_bit_math_h_l1440_c3_43c9_iftrue,
layer6_node0_MUX_bit_math_h_l1440_c3_43c9_iffalse,
layer6_node0_MUX_bit_math_h_l1440_c3_43c9_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 sel,
 in0,
 in1,
 in2,
 in3,
 in4,
 in5,
 in6,
 in7,
 in8,
 in9,
 in10,
 in11,
 in12,
 in13,
 in14,
 in15,
 in16,
 in17,
 in18,
 in19,
 in20,
 in21,
 in22,
 in23,
 in24,
 in25,
 in26,
 in27,
 in28,
 in29,
 in30,
 in31,
 in32,
 in33,
 in34,
 in35,
 in36,
 in37,
 in38,
 in39,
 in40,
 in41,
 in42,
 in43,
 in44,
 in45,
 in46,
 in47,
 in48,
 in49,
 in50,
 in51,
 in52,
 in53,
 in54,
 in55,
 in56,
 in57,
 in58,
 in59,
 in60,
 in61,
 in62,
 in63,
 in64,
 in65,
 in66,
 in67,
 in68,
 in69,
 in70,
 in71,
 in72,
 in73,
 in74,
 in75,
 in76,
 in77,
 in78,
 in79,
 in80,
 in81,
 in82,
 in83,
 in84,
 in85,
 in86,
 in87,
 in88,
 in89,
 in90,
 in91,
 in92,
 in93,
 in94,
 in95,
 in96,
 in97,
 in98,
 in99,
 in100,
 in101,
 in102,
 in103,
 in104,
 in105,
 in106,
 in107,
 in108,
 in109,
 in110,
 in111,
 in112,
 in113,
 in114,
 in115,
 in116,
 in117,
 in118,
 in119,
 in120,
 in121,
 in122,
 in123,
 in124,
 in125,
 in126,
 in127,
 -- All submodule outputs
 layer0_node0_MUX_bit_math_h_l18_c3_ce9b_return_output,
 layer0_node1_MUX_bit_math_h_l29_c3_0e94_return_output,
 layer0_node2_MUX_bit_math_h_l40_c3_e2d9_return_output,
 layer0_node3_MUX_bit_math_h_l51_c3_edc9_return_output,
 layer0_node4_MUX_bit_math_h_l62_c3_f389_return_output,
 layer0_node5_MUX_bit_math_h_l73_c3_d655_return_output,
 layer0_node6_MUX_bit_math_h_l84_c3_5cd3_return_output,
 layer0_node7_MUX_bit_math_h_l95_c3_5030_return_output,
 layer0_node8_MUX_bit_math_h_l106_c3_32cb_return_output,
 layer0_node9_MUX_bit_math_h_l117_c3_4b42_return_output,
 layer0_node10_MUX_bit_math_h_l128_c3_06f3_return_output,
 layer0_node11_MUX_bit_math_h_l139_c3_dbfc_return_output,
 layer0_node12_MUX_bit_math_h_l150_c3_6613_return_output,
 layer0_node13_MUX_bit_math_h_l161_c3_fd42_return_output,
 layer0_node14_MUX_bit_math_h_l172_c3_154a_return_output,
 layer0_node15_MUX_bit_math_h_l183_c3_5274_return_output,
 layer0_node16_MUX_bit_math_h_l194_c3_7a7d_return_output,
 layer0_node17_MUX_bit_math_h_l205_c3_42ac_return_output,
 layer0_node18_MUX_bit_math_h_l216_c3_b8f1_return_output,
 layer0_node19_MUX_bit_math_h_l227_c3_0b12_return_output,
 layer0_node20_MUX_bit_math_h_l238_c3_091e_return_output,
 layer0_node21_MUX_bit_math_h_l249_c3_44d2_return_output,
 layer0_node22_MUX_bit_math_h_l260_c3_db28_return_output,
 layer0_node23_MUX_bit_math_h_l271_c3_0038_return_output,
 layer0_node24_MUX_bit_math_h_l282_c3_1d56_return_output,
 layer0_node25_MUX_bit_math_h_l293_c3_fa3c_return_output,
 layer0_node26_MUX_bit_math_h_l304_c3_220e_return_output,
 layer0_node27_MUX_bit_math_h_l315_c3_37d2_return_output,
 layer0_node28_MUX_bit_math_h_l326_c3_af14_return_output,
 layer0_node29_MUX_bit_math_h_l337_c3_d491_return_output,
 layer0_node30_MUX_bit_math_h_l348_c3_46cf_return_output,
 layer0_node31_MUX_bit_math_h_l359_c3_1ee6_return_output,
 layer0_node32_MUX_bit_math_h_l370_c3_ee39_return_output,
 layer0_node33_MUX_bit_math_h_l381_c3_f57d_return_output,
 layer0_node34_MUX_bit_math_h_l392_c3_8d4e_return_output,
 layer0_node35_MUX_bit_math_h_l403_c3_fa1f_return_output,
 layer0_node36_MUX_bit_math_h_l414_c3_39b4_return_output,
 layer0_node37_MUX_bit_math_h_l425_c3_3900_return_output,
 layer0_node38_MUX_bit_math_h_l436_c3_bea2_return_output,
 layer0_node39_MUX_bit_math_h_l447_c3_3acc_return_output,
 layer0_node40_MUX_bit_math_h_l458_c3_f867_return_output,
 layer0_node41_MUX_bit_math_h_l469_c3_2ffe_return_output,
 layer0_node42_MUX_bit_math_h_l480_c3_1c62_return_output,
 layer0_node43_MUX_bit_math_h_l491_c3_7943_return_output,
 layer0_node44_MUX_bit_math_h_l502_c3_15dc_return_output,
 layer0_node45_MUX_bit_math_h_l513_c3_d638_return_output,
 layer0_node46_MUX_bit_math_h_l524_c3_fdc0_return_output,
 layer0_node47_MUX_bit_math_h_l535_c3_1640_return_output,
 layer0_node48_MUX_bit_math_h_l546_c3_b0f6_return_output,
 layer0_node49_MUX_bit_math_h_l557_c3_adcc_return_output,
 layer0_node50_MUX_bit_math_h_l568_c3_e90e_return_output,
 layer0_node51_MUX_bit_math_h_l579_c3_221f_return_output,
 layer0_node52_MUX_bit_math_h_l590_c3_70e0_return_output,
 layer0_node53_MUX_bit_math_h_l601_c3_e235_return_output,
 layer0_node54_MUX_bit_math_h_l612_c3_f982_return_output,
 layer0_node55_MUX_bit_math_h_l623_c3_bc3d_return_output,
 layer0_node56_MUX_bit_math_h_l634_c3_8e72_return_output,
 layer0_node57_MUX_bit_math_h_l645_c3_0789_return_output,
 layer0_node58_MUX_bit_math_h_l656_c3_d346_return_output,
 layer0_node59_MUX_bit_math_h_l667_c3_d31e_return_output,
 layer0_node60_MUX_bit_math_h_l678_c3_e120_return_output,
 layer0_node61_MUX_bit_math_h_l689_c3_a1a2_return_output,
 layer0_node62_MUX_bit_math_h_l700_c3_4595_return_output,
 layer0_node63_MUX_bit_math_h_l711_c3_c6ab_return_output,
 layer1_node0_MUX_bit_math_h_l728_c3_4268_return_output,
 layer1_node1_MUX_bit_math_h_l739_c3_ff28_return_output,
 layer1_node2_MUX_bit_math_h_l750_c3_543f_return_output,
 layer1_node3_MUX_bit_math_h_l761_c3_5c18_return_output,
 layer1_node4_MUX_bit_math_h_l772_c3_a66b_return_output,
 layer1_node5_MUX_bit_math_h_l783_c3_6db3_return_output,
 layer1_node6_MUX_bit_math_h_l794_c3_4c59_return_output,
 layer1_node7_MUX_bit_math_h_l805_c3_502f_return_output,
 layer1_node8_MUX_bit_math_h_l816_c3_1eec_return_output,
 layer1_node9_MUX_bit_math_h_l827_c3_d105_return_output,
 layer1_node10_MUX_bit_math_h_l838_c3_8a99_return_output,
 layer1_node11_MUX_bit_math_h_l849_c3_e0a5_return_output,
 layer1_node12_MUX_bit_math_h_l860_c3_53b9_return_output,
 layer1_node13_MUX_bit_math_h_l871_c3_672a_return_output,
 layer1_node14_MUX_bit_math_h_l882_c3_2725_return_output,
 layer1_node15_MUX_bit_math_h_l893_c3_b457_return_output,
 layer1_node16_MUX_bit_math_h_l904_c3_8832_return_output,
 layer1_node17_MUX_bit_math_h_l915_c3_0128_return_output,
 layer1_node18_MUX_bit_math_h_l926_c3_a8cf_return_output,
 layer1_node19_MUX_bit_math_h_l937_c3_3d6b_return_output,
 layer1_node20_MUX_bit_math_h_l948_c3_331f_return_output,
 layer1_node21_MUX_bit_math_h_l959_c3_32d5_return_output,
 layer1_node22_MUX_bit_math_h_l970_c3_56f9_return_output,
 layer1_node23_MUX_bit_math_h_l981_c3_251b_return_output,
 layer1_node24_MUX_bit_math_h_l992_c3_a508_return_output,
 layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_return_output,
 layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_return_output,
 layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_return_output,
 layer1_node28_MUX_bit_math_h_l1036_c3_064f_return_output,
 layer1_node29_MUX_bit_math_h_l1047_c3_e950_return_output,
 layer1_node30_MUX_bit_math_h_l1058_c3_fdae_return_output,
 layer1_node31_MUX_bit_math_h_l1069_c3_6030_return_output,
 layer2_node0_MUX_bit_math_h_l1086_c3_122d_return_output,
 layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_return_output,
 layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_return_output,
 layer2_node3_MUX_bit_math_h_l1119_c3_946d_return_output,
 layer2_node4_MUX_bit_math_h_l1130_c3_1f93_return_output,
 layer2_node5_MUX_bit_math_h_l1141_c3_1425_return_output,
 layer2_node6_MUX_bit_math_h_l1152_c3_008a_return_output,
 layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_return_output,
 layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_return_output,
 layer2_node9_MUX_bit_math_h_l1185_c3_98c3_return_output,
 layer2_node10_MUX_bit_math_h_l1196_c3_1666_return_output,
 layer2_node11_MUX_bit_math_h_l1207_c3_b8de_return_output,
 layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_return_output,
 layer2_node13_MUX_bit_math_h_l1229_c3_d585_return_output,
 layer2_node14_MUX_bit_math_h_l1240_c3_beb5_return_output,
 layer2_node15_MUX_bit_math_h_l1251_c3_7550_return_output,
 layer3_node0_MUX_bit_math_h_l1268_c3_302d_return_output,
 layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_return_output,
 layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_return_output,
 layer3_node3_MUX_bit_math_h_l1301_c3_84c3_return_output,
 layer3_node4_MUX_bit_math_h_l1312_c3_8c96_return_output,
 layer3_node5_MUX_bit_math_h_l1323_c3_57ee_return_output,
 layer3_node6_MUX_bit_math_h_l1334_c3_f24c_return_output,
 layer3_node7_MUX_bit_math_h_l1345_c3_c68c_return_output,
 layer4_node0_MUX_bit_math_h_l1362_c3_a122_return_output,
 layer4_node1_MUX_bit_math_h_l1373_c3_c86f_return_output,
 layer4_node2_MUX_bit_math_h_l1384_c3_76f0_return_output,
 layer4_node3_MUX_bit_math_h_l1395_c3_5649_return_output,
 layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_return_output,
 layer5_node1_MUX_bit_math_h_l1423_c3_d92a_return_output,
 layer6_node0_MUX_bit_math_h_l1440_c3_43c9_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(7 downto 0);
 variable VAR_sel : unsigned(6 downto 0);
 variable VAR_in0 : unsigned(7 downto 0);
 variable VAR_in1 : unsigned(7 downto 0);
 variable VAR_in2 : unsigned(7 downto 0);
 variable VAR_in3 : unsigned(7 downto 0);
 variable VAR_in4 : unsigned(7 downto 0);
 variable VAR_in5 : unsigned(7 downto 0);
 variable VAR_in6 : unsigned(7 downto 0);
 variable VAR_in7 : unsigned(7 downto 0);
 variable VAR_in8 : unsigned(7 downto 0);
 variable VAR_in9 : unsigned(7 downto 0);
 variable VAR_in10 : unsigned(7 downto 0);
 variable VAR_in11 : unsigned(7 downto 0);
 variable VAR_in12 : unsigned(7 downto 0);
 variable VAR_in13 : unsigned(7 downto 0);
 variable VAR_in14 : unsigned(7 downto 0);
 variable VAR_in15 : unsigned(7 downto 0);
 variable VAR_in16 : unsigned(7 downto 0);
 variable VAR_in17 : unsigned(7 downto 0);
 variable VAR_in18 : unsigned(7 downto 0);
 variable VAR_in19 : unsigned(7 downto 0);
 variable VAR_in20 : unsigned(7 downto 0);
 variable VAR_in21 : unsigned(7 downto 0);
 variable VAR_in22 : unsigned(7 downto 0);
 variable VAR_in23 : unsigned(7 downto 0);
 variable VAR_in24 : unsigned(7 downto 0);
 variable VAR_in25 : unsigned(7 downto 0);
 variable VAR_in26 : unsigned(7 downto 0);
 variable VAR_in27 : unsigned(7 downto 0);
 variable VAR_in28 : unsigned(7 downto 0);
 variable VAR_in29 : unsigned(7 downto 0);
 variable VAR_in30 : unsigned(7 downto 0);
 variable VAR_in31 : unsigned(7 downto 0);
 variable VAR_in32 : unsigned(7 downto 0);
 variable VAR_in33 : unsigned(7 downto 0);
 variable VAR_in34 : unsigned(7 downto 0);
 variable VAR_in35 : unsigned(7 downto 0);
 variable VAR_in36 : unsigned(7 downto 0);
 variable VAR_in37 : unsigned(7 downto 0);
 variable VAR_in38 : unsigned(7 downto 0);
 variable VAR_in39 : unsigned(7 downto 0);
 variable VAR_in40 : unsigned(7 downto 0);
 variable VAR_in41 : unsigned(7 downto 0);
 variable VAR_in42 : unsigned(7 downto 0);
 variable VAR_in43 : unsigned(7 downto 0);
 variable VAR_in44 : unsigned(7 downto 0);
 variable VAR_in45 : unsigned(7 downto 0);
 variable VAR_in46 : unsigned(7 downto 0);
 variable VAR_in47 : unsigned(7 downto 0);
 variable VAR_in48 : unsigned(7 downto 0);
 variable VAR_in49 : unsigned(7 downto 0);
 variable VAR_in50 : unsigned(7 downto 0);
 variable VAR_in51 : unsigned(7 downto 0);
 variable VAR_in52 : unsigned(7 downto 0);
 variable VAR_in53 : unsigned(7 downto 0);
 variable VAR_in54 : unsigned(7 downto 0);
 variable VAR_in55 : unsigned(7 downto 0);
 variable VAR_in56 : unsigned(7 downto 0);
 variable VAR_in57 : unsigned(7 downto 0);
 variable VAR_in58 : unsigned(7 downto 0);
 variable VAR_in59 : unsigned(7 downto 0);
 variable VAR_in60 : unsigned(7 downto 0);
 variable VAR_in61 : unsigned(7 downto 0);
 variable VAR_in62 : unsigned(7 downto 0);
 variable VAR_in63 : unsigned(7 downto 0);
 variable VAR_in64 : unsigned(7 downto 0);
 variable VAR_in65 : unsigned(7 downto 0);
 variable VAR_in66 : unsigned(7 downto 0);
 variable VAR_in67 : unsigned(7 downto 0);
 variable VAR_in68 : unsigned(7 downto 0);
 variable VAR_in69 : unsigned(7 downto 0);
 variable VAR_in70 : unsigned(7 downto 0);
 variable VAR_in71 : unsigned(7 downto 0);
 variable VAR_in72 : unsigned(7 downto 0);
 variable VAR_in73 : unsigned(7 downto 0);
 variable VAR_in74 : unsigned(7 downto 0);
 variable VAR_in75 : unsigned(7 downto 0);
 variable VAR_in76 : unsigned(7 downto 0);
 variable VAR_in77 : unsigned(7 downto 0);
 variable VAR_in78 : unsigned(7 downto 0);
 variable VAR_in79 : unsigned(7 downto 0);
 variable VAR_in80 : unsigned(7 downto 0);
 variable VAR_in81 : unsigned(7 downto 0);
 variable VAR_in82 : unsigned(7 downto 0);
 variable VAR_in83 : unsigned(7 downto 0);
 variable VAR_in84 : unsigned(7 downto 0);
 variable VAR_in85 : unsigned(7 downto 0);
 variable VAR_in86 : unsigned(7 downto 0);
 variable VAR_in87 : unsigned(7 downto 0);
 variable VAR_in88 : unsigned(7 downto 0);
 variable VAR_in89 : unsigned(7 downto 0);
 variable VAR_in90 : unsigned(7 downto 0);
 variable VAR_in91 : unsigned(7 downto 0);
 variable VAR_in92 : unsigned(7 downto 0);
 variable VAR_in93 : unsigned(7 downto 0);
 variable VAR_in94 : unsigned(7 downto 0);
 variable VAR_in95 : unsigned(7 downto 0);
 variable VAR_in96 : unsigned(7 downto 0);
 variable VAR_in97 : unsigned(7 downto 0);
 variable VAR_in98 : unsigned(7 downto 0);
 variable VAR_in99 : unsigned(7 downto 0);
 variable VAR_in100 : unsigned(7 downto 0);
 variable VAR_in101 : unsigned(7 downto 0);
 variable VAR_in102 : unsigned(7 downto 0);
 variable VAR_in103 : unsigned(7 downto 0);
 variable VAR_in104 : unsigned(7 downto 0);
 variable VAR_in105 : unsigned(7 downto 0);
 variable VAR_in106 : unsigned(7 downto 0);
 variable VAR_in107 : unsigned(7 downto 0);
 variable VAR_in108 : unsigned(7 downto 0);
 variable VAR_in109 : unsigned(7 downto 0);
 variable VAR_in110 : unsigned(7 downto 0);
 variable VAR_in111 : unsigned(7 downto 0);
 variable VAR_in112 : unsigned(7 downto 0);
 variable VAR_in113 : unsigned(7 downto 0);
 variable VAR_in114 : unsigned(7 downto 0);
 variable VAR_in115 : unsigned(7 downto 0);
 variable VAR_in116 : unsigned(7 downto 0);
 variable VAR_in117 : unsigned(7 downto 0);
 variable VAR_in118 : unsigned(7 downto 0);
 variable VAR_in119 : unsigned(7 downto 0);
 variable VAR_in120 : unsigned(7 downto 0);
 variable VAR_in121 : unsigned(7 downto 0);
 variable VAR_in122 : unsigned(7 downto 0);
 variable VAR_in123 : unsigned(7 downto 0);
 variable VAR_in124 : unsigned(7 downto 0);
 variable VAR_in125 : unsigned(7 downto 0);
 variable VAR_in126 : unsigned(7 downto 0);
 variable VAR_in127 : unsigned(7 downto 0);
 variable VAR_sel0 : unsigned(0 downto 0);
 variable VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output : unsigned(0 downto 0);
 variable VAR_layer0_node0 : unsigned(7 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_ce9b_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_ce9b_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_ce9b_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_ce9b_cond : unsigned(0 downto 0);
 variable VAR_layer0_node1 : unsigned(7 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_0e94_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_0e94_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_0e94_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_0e94_cond : unsigned(0 downto 0);
 variable VAR_layer0_node2 : unsigned(7 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_e2d9_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_e2d9_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_e2d9_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_e2d9_cond : unsigned(0 downto 0);
 variable VAR_layer0_node3 : unsigned(7 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_edc9_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_edc9_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_edc9_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_edc9_cond : unsigned(0 downto 0);
 variable VAR_layer0_node4 : unsigned(7 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_f389_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_f389_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_f389_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_f389_cond : unsigned(0 downto 0);
 variable VAR_layer0_node5 : unsigned(7 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_d655_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_d655_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_d655_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_d655_cond : unsigned(0 downto 0);
 variable VAR_layer0_node6 : unsigned(7 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_5cd3_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_5cd3_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_5cd3_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_5cd3_cond : unsigned(0 downto 0);
 variable VAR_layer0_node7 : unsigned(7 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_5030_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_5030_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_5030_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_5030_cond : unsigned(0 downto 0);
 variable VAR_layer0_node8 : unsigned(7 downto 0);
 variable VAR_layer0_node8_MUX_bit_math_h_l106_c3_32cb_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node8_MUX_bit_math_h_l106_c3_32cb_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node8_MUX_bit_math_h_l106_c3_32cb_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node8_MUX_bit_math_h_l106_c3_32cb_cond : unsigned(0 downto 0);
 variable VAR_layer0_node9 : unsigned(7 downto 0);
 variable VAR_layer0_node9_MUX_bit_math_h_l117_c3_4b42_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node9_MUX_bit_math_h_l117_c3_4b42_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node9_MUX_bit_math_h_l117_c3_4b42_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node9_MUX_bit_math_h_l117_c3_4b42_cond : unsigned(0 downto 0);
 variable VAR_layer0_node10 : unsigned(7 downto 0);
 variable VAR_layer0_node10_MUX_bit_math_h_l128_c3_06f3_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node10_MUX_bit_math_h_l128_c3_06f3_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node10_MUX_bit_math_h_l128_c3_06f3_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node10_MUX_bit_math_h_l128_c3_06f3_cond : unsigned(0 downto 0);
 variable VAR_layer0_node11 : unsigned(7 downto 0);
 variable VAR_layer0_node11_MUX_bit_math_h_l139_c3_dbfc_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node11_MUX_bit_math_h_l139_c3_dbfc_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node11_MUX_bit_math_h_l139_c3_dbfc_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node11_MUX_bit_math_h_l139_c3_dbfc_cond : unsigned(0 downto 0);
 variable VAR_layer0_node12 : unsigned(7 downto 0);
 variable VAR_layer0_node12_MUX_bit_math_h_l150_c3_6613_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node12_MUX_bit_math_h_l150_c3_6613_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node12_MUX_bit_math_h_l150_c3_6613_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node12_MUX_bit_math_h_l150_c3_6613_cond : unsigned(0 downto 0);
 variable VAR_layer0_node13 : unsigned(7 downto 0);
 variable VAR_layer0_node13_MUX_bit_math_h_l161_c3_fd42_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node13_MUX_bit_math_h_l161_c3_fd42_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node13_MUX_bit_math_h_l161_c3_fd42_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node13_MUX_bit_math_h_l161_c3_fd42_cond : unsigned(0 downto 0);
 variable VAR_layer0_node14 : unsigned(7 downto 0);
 variable VAR_layer0_node14_MUX_bit_math_h_l172_c3_154a_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node14_MUX_bit_math_h_l172_c3_154a_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node14_MUX_bit_math_h_l172_c3_154a_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node14_MUX_bit_math_h_l172_c3_154a_cond : unsigned(0 downto 0);
 variable VAR_layer0_node15 : unsigned(7 downto 0);
 variable VAR_layer0_node15_MUX_bit_math_h_l183_c3_5274_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node15_MUX_bit_math_h_l183_c3_5274_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node15_MUX_bit_math_h_l183_c3_5274_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node15_MUX_bit_math_h_l183_c3_5274_cond : unsigned(0 downto 0);
 variable VAR_layer0_node16 : unsigned(7 downto 0);
 variable VAR_layer0_node16_MUX_bit_math_h_l194_c3_7a7d_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node16_MUX_bit_math_h_l194_c3_7a7d_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node16_MUX_bit_math_h_l194_c3_7a7d_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node16_MUX_bit_math_h_l194_c3_7a7d_cond : unsigned(0 downto 0);
 variable VAR_layer0_node17 : unsigned(7 downto 0);
 variable VAR_layer0_node17_MUX_bit_math_h_l205_c3_42ac_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node17_MUX_bit_math_h_l205_c3_42ac_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node17_MUX_bit_math_h_l205_c3_42ac_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node17_MUX_bit_math_h_l205_c3_42ac_cond : unsigned(0 downto 0);
 variable VAR_layer0_node18 : unsigned(7 downto 0);
 variable VAR_layer0_node18_MUX_bit_math_h_l216_c3_b8f1_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node18_MUX_bit_math_h_l216_c3_b8f1_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node18_MUX_bit_math_h_l216_c3_b8f1_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node18_MUX_bit_math_h_l216_c3_b8f1_cond : unsigned(0 downto 0);
 variable VAR_layer0_node19 : unsigned(7 downto 0);
 variable VAR_layer0_node19_MUX_bit_math_h_l227_c3_0b12_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node19_MUX_bit_math_h_l227_c3_0b12_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node19_MUX_bit_math_h_l227_c3_0b12_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node19_MUX_bit_math_h_l227_c3_0b12_cond : unsigned(0 downto 0);
 variable VAR_layer0_node20 : unsigned(7 downto 0);
 variable VAR_layer0_node20_MUX_bit_math_h_l238_c3_091e_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node20_MUX_bit_math_h_l238_c3_091e_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node20_MUX_bit_math_h_l238_c3_091e_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node20_MUX_bit_math_h_l238_c3_091e_cond : unsigned(0 downto 0);
 variable VAR_layer0_node21 : unsigned(7 downto 0);
 variable VAR_layer0_node21_MUX_bit_math_h_l249_c3_44d2_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node21_MUX_bit_math_h_l249_c3_44d2_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node21_MUX_bit_math_h_l249_c3_44d2_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node21_MUX_bit_math_h_l249_c3_44d2_cond : unsigned(0 downto 0);
 variable VAR_layer0_node22 : unsigned(7 downto 0);
 variable VAR_layer0_node22_MUX_bit_math_h_l260_c3_db28_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node22_MUX_bit_math_h_l260_c3_db28_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node22_MUX_bit_math_h_l260_c3_db28_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node22_MUX_bit_math_h_l260_c3_db28_cond : unsigned(0 downto 0);
 variable VAR_layer0_node23 : unsigned(7 downto 0);
 variable VAR_layer0_node23_MUX_bit_math_h_l271_c3_0038_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node23_MUX_bit_math_h_l271_c3_0038_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node23_MUX_bit_math_h_l271_c3_0038_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node23_MUX_bit_math_h_l271_c3_0038_cond : unsigned(0 downto 0);
 variable VAR_layer0_node24 : unsigned(7 downto 0);
 variable VAR_layer0_node24_MUX_bit_math_h_l282_c3_1d56_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node24_MUX_bit_math_h_l282_c3_1d56_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node24_MUX_bit_math_h_l282_c3_1d56_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node24_MUX_bit_math_h_l282_c3_1d56_cond : unsigned(0 downto 0);
 variable VAR_layer0_node25 : unsigned(7 downto 0);
 variable VAR_layer0_node25_MUX_bit_math_h_l293_c3_fa3c_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node25_MUX_bit_math_h_l293_c3_fa3c_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node25_MUX_bit_math_h_l293_c3_fa3c_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node25_MUX_bit_math_h_l293_c3_fa3c_cond : unsigned(0 downto 0);
 variable VAR_layer0_node26 : unsigned(7 downto 0);
 variable VAR_layer0_node26_MUX_bit_math_h_l304_c3_220e_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node26_MUX_bit_math_h_l304_c3_220e_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node26_MUX_bit_math_h_l304_c3_220e_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node26_MUX_bit_math_h_l304_c3_220e_cond : unsigned(0 downto 0);
 variable VAR_layer0_node27 : unsigned(7 downto 0);
 variable VAR_layer0_node27_MUX_bit_math_h_l315_c3_37d2_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node27_MUX_bit_math_h_l315_c3_37d2_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node27_MUX_bit_math_h_l315_c3_37d2_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node27_MUX_bit_math_h_l315_c3_37d2_cond : unsigned(0 downto 0);
 variable VAR_layer0_node28 : unsigned(7 downto 0);
 variable VAR_layer0_node28_MUX_bit_math_h_l326_c3_af14_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node28_MUX_bit_math_h_l326_c3_af14_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node28_MUX_bit_math_h_l326_c3_af14_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node28_MUX_bit_math_h_l326_c3_af14_cond : unsigned(0 downto 0);
 variable VAR_layer0_node29 : unsigned(7 downto 0);
 variable VAR_layer0_node29_MUX_bit_math_h_l337_c3_d491_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node29_MUX_bit_math_h_l337_c3_d491_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node29_MUX_bit_math_h_l337_c3_d491_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node29_MUX_bit_math_h_l337_c3_d491_cond : unsigned(0 downto 0);
 variable VAR_layer0_node30 : unsigned(7 downto 0);
 variable VAR_layer0_node30_MUX_bit_math_h_l348_c3_46cf_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node30_MUX_bit_math_h_l348_c3_46cf_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node30_MUX_bit_math_h_l348_c3_46cf_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node30_MUX_bit_math_h_l348_c3_46cf_cond : unsigned(0 downto 0);
 variable VAR_layer0_node31 : unsigned(7 downto 0);
 variable VAR_layer0_node31_MUX_bit_math_h_l359_c3_1ee6_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node31_MUX_bit_math_h_l359_c3_1ee6_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node31_MUX_bit_math_h_l359_c3_1ee6_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node31_MUX_bit_math_h_l359_c3_1ee6_cond : unsigned(0 downto 0);
 variable VAR_layer0_node32 : unsigned(7 downto 0);
 variable VAR_layer0_node32_MUX_bit_math_h_l370_c3_ee39_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node32_MUX_bit_math_h_l370_c3_ee39_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node32_MUX_bit_math_h_l370_c3_ee39_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node32_MUX_bit_math_h_l370_c3_ee39_cond : unsigned(0 downto 0);
 variable VAR_layer0_node33 : unsigned(7 downto 0);
 variable VAR_layer0_node33_MUX_bit_math_h_l381_c3_f57d_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node33_MUX_bit_math_h_l381_c3_f57d_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node33_MUX_bit_math_h_l381_c3_f57d_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node33_MUX_bit_math_h_l381_c3_f57d_cond : unsigned(0 downto 0);
 variable VAR_layer0_node34 : unsigned(7 downto 0);
 variable VAR_layer0_node34_MUX_bit_math_h_l392_c3_8d4e_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node34_MUX_bit_math_h_l392_c3_8d4e_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node34_MUX_bit_math_h_l392_c3_8d4e_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node34_MUX_bit_math_h_l392_c3_8d4e_cond : unsigned(0 downto 0);
 variable VAR_layer0_node35 : unsigned(7 downto 0);
 variable VAR_layer0_node35_MUX_bit_math_h_l403_c3_fa1f_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node35_MUX_bit_math_h_l403_c3_fa1f_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node35_MUX_bit_math_h_l403_c3_fa1f_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node35_MUX_bit_math_h_l403_c3_fa1f_cond : unsigned(0 downto 0);
 variable VAR_layer0_node36 : unsigned(7 downto 0);
 variable VAR_layer0_node36_MUX_bit_math_h_l414_c3_39b4_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node36_MUX_bit_math_h_l414_c3_39b4_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node36_MUX_bit_math_h_l414_c3_39b4_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node36_MUX_bit_math_h_l414_c3_39b4_cond : unsigned(0 downto 0);
 variable VAR_layer0_node37 : unsigned(7 downto 0);
 variable VAR_layer0_node37_MUX_bit_math_h_l425_c3_3900_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node37_MUX_bit_math_h_l425_c3_3900_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node37_MUX_bit_math_h_l425_c3_3900_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node37_MUX_bit_math_h_l425_c3_3900_cond : unsigned(0 downto 0);
 variable VAR_layer0_node38 : unsigned(7 downto 0);
 variable VAR_layer0_node38_MUX_bit_math_h_l436_c3_bea2_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node38_MUX_bit_math_h_l436_c3_bea2_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node38_MUX_bit_math_h_l436_c3_bea2_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node38_MUX_bit_math_h_l436_c3_bea2_cond : unsigned(0 downto 0);
 variable VAR_layer0_node39 : unsigned(7 downto 0);
 variable VAR_layer0_node39_MUX_bit_math_h_l447_c3_3acc_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node39_MUX_bit_math_h_l447_c3_3acc_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node39_MUX_bit_math_h_l447_c3_3acc_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node39_MUX_bit_math_h_l447_c3_3acc_cond : unsigned(0 downto 0);
 variable VAR_layer0_node40 : unsigned(7 downto 0);
 variable VAR_layer0_node40_MUX_bit_math_h_l458_c3_f867_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node40_MUX_bit_math_h_l458_c3_f867_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node40_MUX_bit_math_h_l458_c3_f867_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node40_MUX_bit_math_h_l458_c3_f867_cond : unsigned(0 downto 0);
 variable VAR_layer0_node41 : unsigned(7 downto 0);
 variable VAR_layer0_node41_MUX_bit_math_h_l469_c3_2ffe_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node41_MUX_bit_math_h_l469_c3_2ffe_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node41_MUX_bit_math_h_l469_c3_2ffe_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node41_MUX_bit_math_h_l469_c3_2ffe_cond : unsigned(0 downto 0);
 variable VAR_layer0_node42 : unsigned(7 downto 0);
 variable VAR_layer0_node42_MUX_bit_math_h_l480_c3_1c62_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node42_MUX_bit_math_h_l480_c3_1c62_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node42_MUX_bit_math_h_l480_c3_1c62_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node42_MUX_bit_math_h_l480_c3_1c62_cond : unsigned(0 downto 0);
 variable VAR_layer0_node43 : unsigned(7 downto 0);
 variable VAR_layer0_node43_MUX_bit_math_h_l491_c3_7943_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node43_MUX_bit_math_h_l491_c3_7943_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node43_MUX_bit_math_h_l491_c3_7943_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node43_MUX_bit_math_h_l491_c3_7943_cond : unsigned(0 downto 0);
 variable VAR_layer0_node44 : unsigned(7 downto 0);
 variable VAR_layer0_node44_MUX_bit_math_h_l502_c3_15dc_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node44_MUX_bit_math_h_l502_c3_15dc_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node44_MUX_bit_math_h_l502_c3_15dc_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node44_MUX_bit_math_h_l502_c3_15dc_cond : unsigned(0 downto 0);
 variable VAR_layer0_node45 : unsigned(7 downto 0);
 variable VAR_layer0_node45_MUX_bit_math_h_l513_c3_d638_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node45_MUX_bit_math_h_l513_c3_d638_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node45_MUX_bit_math_h_l513_c3_d638_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node45_MUX_bit_math_h_l513_c3_d638_cond : unsigned(0 downto 0);
 variable VAR_layer0_node46 : unsigned(7 downto 0);
 variable VAR_layer0_node46_MUX_bit_math_h_l524_c3_fdc0_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node46_MUX_bit_math_h_l524_c3_fdc0_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node46_MUX_bit_math_h_l524_c3_fdc0_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node46_MUX_bit_math_h_l524_c3_fdc0_cond : unsigned(0 downto 0);
 variable VAR_layer0_node47 : unsigned(7 downto 0);
 variable VAR_layer0_node47_MUX_bit_math_h_l535_c3_1640_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node47_MUX_bit_math_h_l535_c3_1640_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node47_MUX_bit_math_h_l535_c3_1640_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node47_MUX_bit_math_h_l535_c3_1640_cond : unsigned(0 downto 0);
 variable VAR_layer0_node48 : unsigned(7 downto 0);
 variable VAR_layer0_node48_MUX_bit_math_h_l546_c3_b0f6_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node48_MUX_bit_math_h_l546_c3_b0f6_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node48_MUX_bit_math_h_l546_c3_b0f6_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node48_MUX_bit_math_h_l546_c3_b0f6_cond : unsigned(0 downto 0);
 variable VAR_layer0_node49 : unsigned(7 downto 0);
 variable VAR_layer0_node49_MUX_bit_math_h_l557_c3_adcc_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node49_MUX_bit_math_h_l557_c3_adcc_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node49_MUX_bit_math_h_l557_c3_adcc_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node49_MUX_bit_math_h_l557_c3_adcc_cond : unsigned(0 downto 0);
 variable VAR_layer0_node50 : unsigned(7 downto 0);
 variable VAR_layer0_node50_MUX_bit_math_h_l568_c3_e90e_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node50_MUX_bit_math_h_l568_c3_e90e_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node50_MUX_bit_math_h_l568_c3_e90e_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node50_MUX_bit_math_h_l568_c3_e90e_cond : unsigned(0 downto 0);
 variable VAR_layer0_node51 : unsigned(7 downto 0);
 variable VAR_layer0_node51_MUX_bit_math_h_l579_c3_221f_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node51_MUX_bit_math_h_l579_c3_221f_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node51_MUX_bit_math_h_l579_c3_221f_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node51_MUX_bit_math_h_l579_c3_221f_cond : unsigned(0 downto 0);
 variable VAR_layer0_node52 : unsigned(7 downto 0);
 variable VAR_layer0_node52_MUX_bit_math_h_l590_c3_70e0_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node52_MUX_bit_math_h_l590_c3_70e0_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node52_MUX_bit_math_h_l590_c3_70e0_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node52_MUX_bit_math_h_l590_c3_70e0_cond : unsigned(0 downto 0);
 variable VAR_layer0_node53 : unsigned(7 downto 0);
 variable VAR_layer0_node53_MUX_bit_math_h_l601_c3_e235_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node53_MUX_bit_math_h_l601_c3_e235_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node53_MUX_bit_math_h_l601_c3_e235_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node53_MUX_bit_math_h_l601_c3_e235_cond : unsigned(0 downto 0);
 variable VAR_layer0_node54 : unsigned(7 downto 0);
 variable VAR_layer0_node54_MUX_bit_math_h_l612_c3_f982_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node54_MUX_bit_math_h_l612_c3_f982_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node54_MUX_bit_math_h_l612_c3_f982_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node54_MUX_bit_math_h_l612_c3_f982_cond : unsigned(0 downto 0);
 variable VAR_layer0_node55 : unsigned(7 downto 0);
 variable VAR_layer0_node55_MUX_bit_math_h_l623_c3_bc3d_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node55_MUX_bit_math_h_l623_c3_bc3d_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node55_MUX_bit_math_h_l623_c3_bc3d_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node55_MUX_bit_math_h_l623_c3_bc3d_cond : unsigned(0 downto 0);
 variable VAR_layer0_node56 : unsigned(7 downto 0);
 variable VAR_layer0_node56_MUX_bit_math_h_l634_c3_8e72_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node56_MUX_bit_math_h_l634_c3_8e72_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node56_MUX_bit_math_h_l634_c3_8e72_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node56_MUX_bit_math_h_l634_c3_8e72_cond : unsigned(0 downto 0);
 variable VAR_layer0_node57 : unsigned(7 downto 0);
 variable VAR_layer0_node57_MUX_bit_math_h_l645_c3_0789_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node57_MUX_bit_math_h_l645_c3_0789_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node57_MUX_bit_math_h_l645_c3_0789_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node57_MUX_bit_math_h_l645_c3_0789_cond : unsigned(0 downto 0);
 variable VAR_layer0_node58 : unsigned(7 downto 0);
 variable VAR_layer0_node58_MUX_bit_math_h_l656_c3_d346_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node58_MUX_bit_math_h_l656_c3_d346_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node58_MUX_bit_math_h_l656_c3_d346_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node58_MUX_bit_math_h_l656_c3_d346_cond : unsigned(0 downto 0);
 variable VAR_layer0_node59 : unsigned(7 downto 0);
 variable VAR_layer0_node59_MUX_bit_math_h_l667_c3_d31e_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node59_MUX_bit_math_h_l667_c3_d31e_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node59_MUX_bit_math_h_l667_c3_d31e_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node59_MUX_bit_math_h_l667_c3_d31e_cond : unsigned(0 downto 0);
 variable VAR_layer0_node60 : unsigned(7 downto 0);
 variable VAR_layer0_node60_MUX_bit_math_h_l678_c3_e120_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node60_MUX_bit_math_h_l678_c3_e120_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node60_MUX_bit_math_h_l678_c3_e120_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node60_MUX_bit_math_h_l678_c3_e120_cond : unsigned(0 downto 0);
 variable VAR_layer0_node61 : unsigned(7 downto 0);
 variable VAR_layer0_node61_MUX_bit_math_h_l689_c3_a1a2_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node61_MUX_bit_math_h_l689_c3_a1a2_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node61_MUX_bit_math_h_l689_c3_a1a2_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node61_MUX_bit_math_h_l689_c3_a1a2_cond : unsigned(0 downto 0);
 variable VAR_layer0_node62 : unsigned(7 downto 0);
 variable VAR_layer0_node62_MUX_bit_math_h_l700_c3_4595_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node62_MUX_bit_math_h_l700_c3_4595_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node62_MUX_bit_math_h_l700_c3_4595_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node62_MUX_bit_math_h_l700_c3_4595_cond : unsigned(0 downto 0);
 variable VAR_layer0_node63 : unsigned(7 downto 0);
 variable VAR_layer0_node63_MUX_bit_math_h_l711_c3_c6ab_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node63_MUX_bit_math_h_l711_c3_c6ab_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node63_MUX_bit_math_h_l711_c3_c6ab_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node63_MUX_bit_math_h_l711_c3_c6ab_cond : unsigned(0 downto 0);
 variable VAR_sel1 : unsigned(0 downto 0);
 variable VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output : unsigned(0 downto 0);
 variable VAR_layer1_node0 : unsigned(7 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l728_c3_4268_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l728_c3_4268_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l728_c3_4268_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l728_c3_4268_cond : unsigned(0 downto 0);
 variable VAR_layer1_node1 : unsigned(7 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l739_c3_ff28_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l739_c3_ff28_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l739_c3_ff28_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l739_c3_ff28_cond : unsigned(0 downto 0);
 variable VAR_layer1_node2 : unsigned(7 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l750_c3_543f_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l750_c3_543f_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l750_c3_543f_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l750_c3_543f_cond : unsigned(0 downto 0);
 variable VAR_layer1_node3 : unsigned(7 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l761_c3_5c18_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l761_c3_5c18_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l761_c3_5c18_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l761_c3_5c18_cond : unsigned(0 downto 0);
 variable VAR_layer1_node4 : unsigned(7 downto 0);
 variable VAR_layer1_node4_MUX_bit_math_h_l772_c3_a66b_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node4_MUX_bit_math_h_l772_c3_a66b_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node4_MUX_bit_math_h_l772_c3_a66b_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node4_MUX_bit_math_h_l772_c3_a66b_cond : unsigned(0 downto 0);
 variable VAR_layer1_node5 : unsigned(7 downto 0);
 variable VAR_layer1_node5_MUX_bit_math_h_l783_c3_6db3_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node5_MUX_bit_math_h_l783_c3_6db3_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node5_MUX_bit_math_h_l783_c3_6db3_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node5_MUX_bit_math_h_l783_c3_6db3_cond : unsigned(0 downto 0);
 variable VAR_layer1_node6 : unsigned(7 downto 0);
 variable VAR_layer1_node6_MUX_bit_math_h_l794_c3_4c59_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node6_MUX_bit_math_h_l794_c3_4c59_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node6_MUX_bit_math_h_l794_c3_4c59_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node6_MUX_bit_math_h_l794_c3_4c59_cond : unsigned(0 downto 0);
 variable VAR_layer1_node7 : unsigned(7 downto 0);
 variable VAR_layer1_node7_MUX_bit_math_h_l805_c3_502f_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node7_MUX_bit_math_h_l805_c3_502f_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node7_MUX_bit_math_h_l805_c3_502f_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node7_MUX_bit_math_h_l805_c3_502f_cond : unsigned(0 downto 0);
 variable VAR_layer1_node8 : unsigned(7 downto 0);
 variable VAR_layer1_node8_MUX_bit_math_h_l816_c3_1eec_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node8_MUX_bit_math_h_l816_c3_1eec_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node8_MUX_bit_math_h_l816_c3_1eec_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node8_MUX_bit_math_h_l816_c3_1eec_cond : unsigned(0 downto 0);
 variable VAR_layer1_node9 : unsigned(7 downto 0);
 variable VAR_layer1_node9_MUX_bit_math_h_l827_c3_d105_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node9_MUX_bit_math_h_l827_c3_d105_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node9_MUX_bit_math_h_l827_c3_d105_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node9_MUX_bit_math_h_l827_c3_d105_cond : unsigned(0 downto 0);
 variable VAR_layer1_node10 : unsigned(7 downto 0);
 variable VAR_layer1_node10_MUX_bit_math_h_l838_c3_8a99_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node10_MUX_bit_math_h_l838_c3_8a99_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node10_MUX_bit_math_h_l838_c3_8a99_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node10_MUX_bit_math_h_l838_c3_8a99_cond : unsigned(0 downto 0);
 variable VAR_layer1_node11 : unsigned(7 downto 0);
 variable VAR_layer1_node11_MUX_bit_math_h_l849_c3_e0a5_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node11_MUX_bit_math_h_l849_c3_e0a5_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node11_MUX_bit_math_h_l849_c3_e0a5_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node11_MUX_bit_math_h_l849_c3_e0a5_cond : unsigned(0 downto 0);
 variable VAR_layer1_node12 : unsigned(7 downto 0);
 variable VAR_layer1_node12_MUX_bit_math_h_l860_c3_53b9_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node12_MUX_bit_math_h_l860_c3_53b9_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node12_MUX_bit_math_h_l860_c3_53b9_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node12_MUX_bit_math_h_l860_c3_53b9_cond : unsigned(0 downto 0);
 variable VAR_layer1_node13 : unsigned(7 downto 0);
 variable VAR_layer1_node13_MUX_bit_math_h_l871_c3_672a_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node13_MUX_bit_math_h_l871_c3_672a_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node13_MUX_bit_math_h_l871_c3_672a_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node13_MUX_bit_math_h_l871_c3_672a_cond : unsigned(0 downto 0);
 variable VAR_layer1_node14 : unsigned(7 downto 0);
 variable VAR_layer1_node14_MUX_bit_math_h_l882_c3_2725_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node14_MUX_bit_math_h_l882_c3_2725_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node14_MUX_bit_math_h_l882_c3_2725_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node14_MUX_bit_math_h_l882_c3_2725_cond : unsigned(0 downto 0);
 variable VAR_layer1_node15 : unsigned(7 downto 0);
 variable VAR_layer1_node15_MUX_bit_math_h_l893_c3_b457_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node15_MUX_bit_math_h_l893_c3_b457_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node15_MUX_bit_math_h_l893_c3_b457_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node15_MUX_bit_math_h_l893_c3_b457_cond : unsigned(0 downto 0);
 variable VAR_layer1_node16 : unsigned(7 downto 0);
 variable VAR_layer1_node16_MUX_bit_math_h_l904_c3_8832_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node16_MUX_bit_math_h_l904_c3_8832_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node16_MUX_bit_math_h_l904_c3_8832_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node16_MUX_bit_math_h_l904_c3_8832_cond : unsigned(0 downto 0);
 variable VAR_layer1_node17 : unsigned(7 downto 0);
 variable VAR_layer1_node17_MUX_bit_math_h_l915_c3_0128_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node17_MUX_bit_math_h_l915_c3_0128_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node17_MUX_bit_math_h_l915_c3_0128_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node17_MUX_bit_math_h_l915_c3_0128_cond : unsigned(0 downto 0);
 variable VAR_layer1_node18 : unsigned(7 downto 0);
 variable VAR_layer1_node18_MUX_bit_math_h_l926_c3_a8cf_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node18_MUX_bit_math_h_l926_c3_a8cf_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node18_MUX_bit_math_h_l926_c3_a8cf_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node18_MUX_bit_math_h_l926_c3_a8cf_cond : unsigned(0 downto 0);
 variable VAR_layer1_node19 : unsigned(7 downto 0);
 variable VAR_layer1_node19_MUX_bit_math_h_l937_c3_3d6b_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node19_MUX_bit_math_h_l937_c3_3d6b_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node19_MUX_bit_math_h_l937_c3_3d6b_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node19_MUX_bit_math_h_l937_c3_3d6b_cond : unsigned(0 downto 0);
 variable VAR_layer1_node20 : unsigned(7 downto 0);
 variable VAR_layer1_node20_MUX_bit_math_h_l948_c3_331f_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node20_MUX_bit_math_h_l948_c3_331f_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node20_MUX_bit_math_h_l948_c3_331f_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node20_MUX_bit_math_h_l948_c3_331f_cond : unsigned(0 downto 0);
 variable VAR_layer1_node21 : unsigned(7 downto 0);
 variable VAR_layer1_node21_MUX_bit_math_h_l959_c3_32d5_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node21_MUX_bit_math_h_l959_c3_32d5_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node21_MUX_bit_math_h_l959_c3_32d5_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node21_MUX_bit_math_h_l959_c3_32d5_cond : unsigned(0 downto 0);
 variable VAR_layer1_node22 : unsigned(7 downto 0);
 variable VAR_layer1_node22_MUX_bit_math_h_l970_c3_56f9_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node22_MUX_bit_math_h_l970_c3_56f9_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node22_MUX_bit_math_h_l970_c3_56f9_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node22_MUX_bit_math_h_l970_c3_56f9_cond : unsigned(0 downto 0);
 variable VAR_layer1_node23 : unsigned(7 downto 0);
 variable VAR_layer1_node23_MUX_bit_math_h_l981_c3_251b_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node23_MUX_bit_math_h_l981_c3_251b_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node23_MUX_bit_math_h_l981_c3_251b_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node23_MUX_bit_math_h_l981_c3_251b_cond : unsigned(0 downto 0);
 variable VAR_layer1_node24 : unsigned(7 downto 0);
 variable VAR_layer1_node24_MUX_bit_math_h_l992_c3_a508_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node24_MUX_bit_math_h_l992_c3_a508_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node24_MUX_bit_math_h_l992_c3_a508_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node24_MUX_bit_math_h_l992_c3_a508_cond : unsigned(0 downto 0);
 variable VAR_layer1_node25 : unsigned(7 downto 0);
 variable VAR_layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_cond : unsigned(0 downto 0);
 variable VAR_layer1_node26 : unsigned(7 downto 0);
 variable VAR_layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_cond : unsigned(0 downto 0);
 variable VAR_layer1_node27 : unsigned(7 downto 0);
 variable VAR_layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_cond : unsigned(0 downto 0);
 variable VAR_layer1_node28 : unsigned(7 downto 0);
 variable VAR_layer1_node28_MUX_bit_math_h_l1036_c3_064f_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node28_MUX_bit_math_h_l1036_c3_064f_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node28_MUX_bit_math_h_l1036_c3_064f_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node28_MUX_bit_math_h_l1036_c3_064f_cond : unsigned(0 downto 0);
 variable VAR_layer1_node29 : unsigned(7 downto 0);
 variable VAR_layer1_node29_MUX_bit_math_h_l1047_c3_e950_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node29_MUX_bit_math_h_l1047_c3_e950_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node29_MUX_bit_math_h_l1047_c3_e950_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node29_MUX_bit_math_h_l1047_c3_e950_cond : unsigned(0 downto 0);
 variable VAR_layer1_node30 : unsigned(7 downto 0);
 variable VAR_layer1_node30_MUX_bit_math_h_l1058_c3_fdae_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node30_MUX_bit_math_h_l1058_c3_fdae_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node30_MUX_bit_math_h_l1058_c3_fdae_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node30_MUX_bit_math_h_l1058_c3_fdae_cond : unsigned(0 downto 0);
 variable VAR_layer1_node31 : unsigned(7 downto 0);
 variable VAR_layer1_node31_MUX_bit_math_h_l1069_c3_6030_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node31_MUX_bit_math_h_l1069_c3_6030_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node31_MUX_bit_math_h_l1069_c3_6030_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node31_MUX_bit_math_h_l1069_c3_6030_cond : unsigned(0 downto 0);
 variable VAR_sel2 : unsigned(0 downto 0);
 variable VAR_uint7_2_2_bit_math_h_l1082_c10_87dc_return_output : unsigned(0 downto 0);
 variable VAR_layer2_node0 : unsigned(7 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l1086_c3_122d_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l1086_c3_122d_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l1086_c3_122d_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l1086_c3_122d_cond : unsigned(0 downto 0);
 variable VAR_layer2_node1 : unsigned(7 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_cond : unsigned(0 downto 0);
 variable VAR_layer2_node2 : unsigned(7 downto 0);
 variable VAR_layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_cond : unsigned(0 downto 0);
 variable VAR_layer2_node3 : unsigned(7 downto 0);
 variable VAR_layer2_node3_MUX_bit_math_h_l1119_c3_946d_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node3_MUX_bit_math_h_l1119_c3_946d_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node3_MUX_bit_math_h_l1119_c3_946d_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node3_MUX_bit_math_h_l1119_c3_946d_cond : unsigned(0 downto 0);
 variable VAR_layer2_node4 : unsigned(7 downto 0);
 variable VAR_layer2_node4_MUX_bit_math_h_l1130_c3_1f93_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node4_MUX_bit_math_h_l1130_c3_1f93_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node4_MUX_bit_math_h_l1130_c3_1f93_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node4_MUX_bit_math_h_l1130_c3_1f93_cond : unsigned(0 downto 0);
 variable VAR_layer2_node5 : unsigned(7 downto 0);
 variable VAR_layer2_node5_MUX_bit_math_h_l1141_c3_1425_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node5_MUX_bit_math_h_l1141_c3_1425_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node5_MUX_bit_math_h_l1141_c3_1425_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node5_MUX_bit_math_h_l1141_c3_1425_cond : unsigned(0 downto 0);
 variable VAR_layer2_node6 : unsigned(7 downto 0);
 variable VAR_layer2_node6_MUX_bit_math_h_l1152_c3_008a_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node6_MUX_bit_math_h_l1152_c3_008a_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node6_MUX_bit_math_h_l1152_c3_008a_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node6_MUX_bit_math_h_l1152_c3_008a_cond : unsigned(0 downto 0);
 variable VAR_layer2_node7 : unsigned(7 downto 0);
 variable VAR_layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_cond : unsigned(0 downto 0);
 variable VAR_layer2_node8 : unsigned(7 downto 0);
 variable VAR_layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_cond : unsigned(0 downto 0);
 variable VAR_layer2_node9 : unsigned(7 downto 0);
 variable VAR_layer2_node9_MUX_bit_math_h_l1185_c3_98c3_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node9_MUX_bit_math_h_l1185_c3_98c3_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node9_MUX_bit_math_h_l1185_c3_98c3_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node9_MUX_bit_math_h_l1185_c3_98c3_cond : unsigned(0 downto 0);
 variable VAR_layer2_node10 : unsigned(7 downto 0);
 variable VAR_layer2_node10_MUX_bit_math_h_l1196_c3_1666_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node10_MUX_bit_math_h_l1196_c3_1666_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node10_MUX_bit_math_h_l1196_c3_1666_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node10_MUX_bit_math_h_l1196_c3_1666_cond : unsigned(0 downto 0);
 variable VAR_layer2_node11 : unsigned(7 downto 0);
 variable VAR_layer2_node11_MUX_bit_math_h_l1207_c3_b8de_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node11_MUX_bit_math_h_l1207_c3_b8de_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node11_MUX_bit_math_h_l1207_c3_b8de_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node11_MUX_bit_math_h_l1207_c3_b8de_cond : unsigned(0 downto 0);
 variable VAR_layer2_node12 : unsigned(7 downto 0);
 variable VAR_layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_cond : unsigned(0 downto 0);
 variable VAR_layer2_node13 : unsigned(7 downto 0);
 variable VAR_layer2_node13_MUX_bit_math_h_l1229_c3_d585_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node13_MUX_bit_math_h_l1229_c3_d585_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node13_MUX_bit_math_h_l1229_c3_d585_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node13_MUX_bit_math_h_l1229_c3_d585_cond : unsigned(0 downto 0);
 variable VAR_layer2_node14 : unsigned(7 downto 0);
 variable VAR_layer2_node14_MUX_bit_math_h_l1240_c3_beb5_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node14_MUX_bit_math_h_l1240_c3_beb5_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node14_MUX_bit_math_h_l1240_c3_beb5_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node14_MUX_bit_math_h_l1240_c3_beb5_cond : unsigned(0 downto 0);
 variable VAR_layer2_node15 : unsigned(7 downto 0);
 variable VAR_layer2_node15_MUX_bit_math_h_l1251_c3_7550_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node15_MUX_bit_math_h_l1251_c3_7550_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node15_MUX_bit_math_h_l1251_c3_7550_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node15_MUX_bit_math_h_l1251_c3_7550_cond : unsigned(0 downto 0);
 variable VAR_sel3 : unsigned(0 downto 0);
 variable VAR_uint7_3_3_bit_math_h_l1264_c10_51ff_return_output : unsigned(0 downto 0);
 variable VAR_layer3_node0 : unsigned(7 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l1268_c3_302d_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l1268_c3_302d_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l1268_c3_302d_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l1268_c3_302d_cond : unsigned(0 downto 0);
 variable VAR_layer3_node1 : unsigned(7 downto 0);
 variable VAR_layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_cond : unsigned(0 downto 0);
 variable VAR_layer3_node2 : unsigned(7 downto 0);
 variable VAR_layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_cond : unsigned(0 downto 0);
 variable VAR_layer3_node3 : unsigned(7 downto 0);
 variable VAR_layer3_node3_MUX_bit_math_h_l1301_c3_84c3_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node3_MUX_bit_math_h_l1301_c3_84c3_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node3_MUX_bit_math_h_l1301_c3_84c3_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node3_MUX_bit_math_h_l1301_c3_84c3_cond : unsigned(0 downto 0);
 variable VAR_layer3_node4 : unsigned(7 downto 0);
 variable VAR_layer3_node4_MUX_bit_math_h_l1312_c3_8c96_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node4_MUX_bit_math_h_l1312_c3_8c96_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node4_MUX_bit_math_h_l1312_c3_8c96_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node4_MUX_bit_math_h_l1312_c3_8c96_cond : unsigned(0 downto 0);
 variable VAR_layer3_node5 : unsigned(7 downto 0);
 variable VAR_layer3_node5_MUX_bit_math_h_l1323_c3_57ee_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node5_MUX_bit_math_h_l1323_c3_57ee_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node5_MUX_bit_math_h_l1323_c3_57ee_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node5_MUX_bit_math_h_l1323_c3_57ee_cond : unsigned(0 downto 0);
 variable VAR_layer3_node6 : unsigned(7 downto 0);
 variable VAR_layer3_node6_MUX_bit_math_h_l1334_c3_f24c_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node6_MUX_bit_math_h_l1334_c3_f24c_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node6_MUX_bit_math_h_l1334_c3_f24c_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node6_MUX_bit_math_h_l1334_c3_f24c_cond : unsigned(0 downto 0);
 variable VAR_layer3_node7 : unsigned(7 downto 0);
 variable VAR_layer3_node7_MUX_bit_math_h_l1345_c3_c68c_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node7_MUX_bit_math_h_l1345_c3_c68c_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node7_MUX_bit_math_h_l1345_c3_c68c_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node7_MUX_bit_math_h_l1345_c3_c68c_cond : unsigned(0 downto 0);
 variable VAR_sel4 : unsigned(0 downto 0);
 variable VAR_uint7_4_4_bit_math_h_l1358_c10_29af_return_output : unsigned(0 downto 0);
 variable VAR_layer4_node0 : unsigned(7 downto 0);
 variable VAR_layer4_node0_MUX_bit_math_h_l1362_c3_a122_iftrue : unsigned(7 downto 0);
 variable VAR_layer4_node0_MUX_bit_math_h_l1362_c3_a122_iffalse : unsigned(7 downto 0);
 variable VAR_layer4_node0_MUX_bit_math_h_l1362_c3_a122_return_output : unsigned(7 downto 0);
 variable VAR_layer4_node0_MUX_bit_math_h_l1362_c3_a122_cond : unsigned(0 downto 0);
 variable VAR_layer4_node1 : unsigned(7 downto 0);
 variable VAR_layer4_node1_MUX_bit_math_h_l1373_c3_c86f_iftrue : unsigned(7 downto 0);
 variable VAR_layer4_node1_MUX_bit_math_h_l1373_c3_c86f_iffalse : unsigned(7 downto 0);
 variable VAR_layer4_node1_MUX_bit_math_h_l1373_c3_c86f_return_output : unsigned(7 downto 0);
 variable VAR_layer4_node1_MUX_bit_math_h_l1373_c3_c86f_cond : unsigned(0 downto 0);
 variable VAR_layer4_node2 : unsigned(7 downto 0);
 variable VAR_layer4_node2_MUX_bit_math_h_l1384_c3_76f0_iftrue : unsigned(7 downto 0);
 variable VAR_layer4_node2_MUX_bit_math_h_l1384_c3_76f0_iffalse : unsigned(7 downto 0);
 variable VAR_layer4_node2_MUX_bit_math_h_l1384_c3_76f0_return_output : unsigned(7 downto 0);
 variable VAR_layer4_node2_MUX_bit_math_h_l1384_c3_76f0_cond : unsigned(0 downto 0);
 variable VAR_layer4_node3 : unsigned(7 downto 0);
 variable VAR_layer4_node3_MUX_bit_math_h_l1395_c3_5649_iftrue : unsigned(7 downto 0);
 variable VAR_layer4_node3_MUX_bit_math_h_l1395_c3_5649_iffalse : unsigned(7 downto 0);
 variable VAR_layer4_node3_MUX_bit_math_h_l1395_c3_5649_return_output : unsigned(7 downto 0);
 variable VAR_layer4_node3_MUX_bit_math_h_l1395_c3_5649_cond : unsigned(0 downto 0);
 variable VAR_sel5 : unsigned(0 downto 0);
 variable VAR_uint7_5_5_bit_math_h_l1408_c10_a313_return_output : unsigned(0 downto 0);
 variable VAR_layer5_node0 : unsigned(7 downto 0);
 variable VAR_layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_iftrue : unsigned(7 downto 0);
 variable VAR_layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_iffalse : unsigned(7 downto 0);
 variable VAR_layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_return_output : unsigned(7 downto 0);
 variable VAR_layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_cond : unsigned(0 downto 0);
 variable VAR_layer5_node1 : unsigned(7 downto 0);
 variable VAR_layer5_node1_MUX_bit_math_h_l1423_c3_d92a_iftrue : unsigned(7 downto 0);
 variable VAR_layer5_node1_MUX_bit_math_h_l1423_c3_d92a_iffalse : unsigned(7 downto 0);
 variable VAR_layer5_node1_MUX_bit_math_h_l1423_c3_d92a_return_output : unsigned(7 downto 0);
 variable VAR_layer5_node1_MUX_bit_math_h_l1423_c3_d92a_cond : unsigned(0 downto 0);
 variable VAR_sel6 : unsigned(0 downto 0);
 variable VAR_uint7_6_6_bit_math_h_l1436_c10_2ac3_return_output : unsigned(0 downto 0);
 variable VAR_layer6_node0 : unsigned(7 downto 0);
 variable VAR_layer6_node0_MUX_bit_math_h_l1440_c3_43c9_iftrue : unsigned(7 downto 0);
 variable VAR_layer6_node0_MUX_bit_math_h_l1440_c3_43c9_iffalse : unsigned(7 downto 0);
 variable VAR_layer6_node0_MUX_bit_math_h_l1440_c3_43c9_return_output : unsigned(7 downto 0);
 variable VAR_layer6_node0_MUX_bit_math_h_l1440_c3_43c9_cond : unsigned(0 downto 0);
begin

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_sel := sel;
     VAR_in0 := in0;
     VAR_in1 := in1;
     VAR_in2 := in2;
     VAR_in3 := in3;
     VAR_in4 := in4;
     VAR_in5 := in5;
     VAR_in6 := in6;
     VAR_in7 := in7;
     VAR_in8 := in8;
     VAR_in9 := in9;
     VAR_in10 := in10;
     VAR_in11 := in11;
     VAR_in12 := in12;
     VAR_in13 := in13;
     VAR_in14 := in14;
     VAR_in15 := in15;
     VAR_in16 := in16;
     VAR_in17 := in17;
     VAR_in18 := in18;
     VAR_in19 := in19;
     VAR_in20 := in20;
     VAR_in21 := in21;
     VAR_in22 := in22;
     VAR_in23 := in23;
     VAR_in24 := in24;
     VAR_in25 := in25;
     VAR_in26 := in26;
     VAR_in27 := in27;
     VAR_in28 := in28;
     VAR_in29 := in29;
     VAR_in30 := in30;
     VAR_in31 := in31;
     VAR_in32 := in32;
     VAR_in33 := in33;
     VAR_in34 := in34;
     VAR_in35 := in35;
     VAR_in36 := in36;
     VAR_in37 := in37;
     VAR_in38 := in38;
     VAR_in39 := in39;
     VAR_in40 := in40;
     VAR_in41 := in41;
     VAR_in42 := in42;
     VAR_in43 := in43;
     VAR_in44 := in44;
     VAR_in45 := in45;
     VAR_in46 := in46;
     VAR_in47 := in47;
     VAR_in48 := in48;
     VAR_in49 := in49;
     VAR_in50 := in50;
     VAR_in51 := in51;
     VAR_in52 := in52;
     VAR_in53 := in53;
     VAR_in54 := in54;
     VAR_in55 := in55;
     VAR_in56 := in56;
     VAR_in57 := in57;
     VAR_in58 := in58;
     VAR_in59 := in59;
     VAR_in60 := in60;
     VAR_in61 := in61;
     VAR_in62 := in62;
     VAR_in63 := in63;
     VAR_in64 := in64;
     VAR_in65 := in65;
     VAR_in66 := in66;
     VAR_in67 := in67;
     VAR_in68 := in68;
     VAR_in69 := in69;
     VAR_in70 := in70;
     VAR_in71 := in71;
     VAR_in72 := in72;
     VAR_in73 := in73;
     VAR_in74 := in74;
     VAR_in75 := in75;
     VAR_in76 := in76;
     VAR_in77 := in77;
     VAR_in78 := in78;
     VAR_in79 := in79;
     VAR_in80 := in80;
     VAR_in81 := in81;
     VAR_in82 := in82;
     VAR_in83 := in83;
     VAR_in84 := in84;
     VAR_in85 := in85;
     VAR_in86 := in86;
     VAR_in87 := in87;
     VAR_in88 := in88;
     VAR_in89 := in89;
     VAR_in90 := in90;
     VAR_in91 := in91;
     VAR_in92 := in92;
     VAR_in93 := in93;
     VAR_in94 := in94;
     VAR_in95 := in95;
     VAR_in96 := in96;
     VAR_in97 := in97;
     VAR_in98 := in98;
     VAR_in99 := in99;
     VAR_in100 := in100;
     VAR_in101 := in101;
     VAR_in102 := in102;
     VAR_in103 := in103;
     VAR_in104 := in104;
     VAR_in105 := in105;
     VAR_in106 := in106;
     VAR_in107 := in107;
     VAR_in108 := in108;
     VAR_in109 := in109;
     VAR_in110 := in110;
     VAR_in111 := in111;
     VAR_in112 := in112;
     VAR_in113 := in113;
     VAR_in114 := in114;
     VAR_in115 := in115;
     VAR_in116 := in116;
     VAR_in117 := in117;
     VAR_in118 := in118;
     VAR_in119 := in119;
     VAR_in120 := in120;
     VAR_in121 := in121;
     VAR_in122 := in122;
     VAR_in123 := in123;
     VAR_in124 := in124;
     VAR_in125 := in125;
     VAR_in126 := in126;
     VAR_in127 := in127;

     -- Submodule level 0
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_ce9b_iffalse := VAR_in0;
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_ce9b_iftrue := VAR_in1;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_d655_iffalse := VAR_in10;
     VAR_layer0_node50_MUX_bit_math_h_l568_c3_e90e_iffalse := VAR_in100;
     VAR_layer0_node50_MUX_bit_math_h_l568_c3_e90e_iftrue := VAR_in101;
     VAR_layer0_node51_MUX_bit_math_h_l579_c3_221f_iffalse := VAR_in102;
     VAR_layer0_node51_MUX_bit_math_h_l579_c3_221f_iftrue := VAR_in103;
     VAR_layer0_node52_MUX_bit_math_h_l590_c3_70e0_iffalse := VAR_in104;
     VAR_layer0_node52_MUX_bit_math_h_l590_c3_70e0_iftrue := VAR_in105;
     VAR_layer0_node53_MUX_bit_math_h_l601_c3_e235_iffalse := VAR_in106;
     VAR_layer0_node53_MUX_bit_math_h_l601_c3_e235_iftrue := VAR_in107;
     VAR_layer0_node54_MUX_bit_math_h_l612_c3_f982_iffalse := VAR_in108;
     VAR_layer0_node54_MUX_bit_math_h_l612_c3_f982_iftrue := VAR_in109;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_d655_iftrue := VAR_in11;
     VAR_layer0_node55_MUX_bit_math_h_l623_c3_bc3d_iffalse := VAR_in110;
     VAR_layer0_node55_MUX_bit_math_h_l623_c3_bc3d_iftrue := VAR_in111;
     VAR_layer0_node56_MUX_bit_math_h_l634_c3_8e72_iffalse := VAR_in112;
     VAR_layer0_node56_MUX_bit_math_h_l634_c3_8e72_iftrue := VAR_in113;
     VAR_layer0_node57_MUX_bit_math_h_l645_c3_0789_iffalse := VAR_in114;
     VAR_layer0_node57_MUX_bit_math_h_l645_c3_0789_iftrue := VAR_in115;
     VAR_layer0_node58_MUX_bit_math_h_l656_c3_d346_iffalse := VAR_in116;
     VAR_layer0_node58_MUX_bit_math_h_l656_c3_d346_iftrue := VAR_in117;
     VAR_layer0_node59_MUX_bit_math_h_l667_c3_d31e_iffalse := VAR_in118;
     VAR_layer0_node59_MUX_bit_math_h_l667_c3_d31e_iftrue := VAR_in119;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_5cd3_iffalse := VAR_in12;
     VAR_layer0_node60_MUX_bit_math_h_l678_c3_e120_iffalse := VAR_in120;
     VAR_layer0_node60_MUX_bit_math_h_l678_c3_e120_iftrue := VAR_in121;
     VAR_layer0_node61_MUX_bit_math_h_l689_c3_a1a2_iffalse := VAR_in122;
     VAR_layer0_node61_MUX_bit_math_h_l689_c3_a1a2_iftrue := VAR_in123;
     VAR_layer0_node62_MUX_bit_math_h_l700_c3_4595_iffalse := VAR_in124;
     VAR_layer0_node62_MUX_bit_math_h_l700_c3_4595_iftrue := VAR_in125;
     VAR_layer0_node63_MUX_bit_math_h_l711_c3_c6ab_iffalse := VAR_in126;
     VAR_layer0_node63_MUX_bit_math_h_l711_c3_c6ab_iftrue := VAR_in127;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_5cd3_iftrue := VAR_in13;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_5030_iffalse := VAR_in14;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_5030_iftrue := VAR_in15;
     VAR_layer0_node8_MUX_bit_math_h_l106_c3_32cb_iffalse := VAR_in16;
     VAR_layer0_node8_MUX_bit_math_h_l106_c3_32cb_iftrue := VAR_in17;
     VAR_layer0_node9_MUX_bit_math_h_l117_c3_4b42_iffalse := VAR_in18;
     VAR_layer0_node9_MUX_bit_math_h_l117_c3_4b42_iftrue := VAR_in19;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_0e94_iffalse := VAR_in2;
     VAR_layer0_node10_MUX_bit_math_h_l128_c3_06f3_iffalse := VAR_in20;
     VAR_layer0_node10_MUX_bit_math_h_l128_c3_06f3_iftrue := VAR_in21;
     VAR_layer0_node11_MUX_bit_math_h_l139_c3_dbfc_iffalse := VAR_in22;
     VAR_layer0_node11_MUX_bit_math_h_l139_c3_dbfc_iftrue := VAR_in23;
     VAR_layer0_node12_MUX_bit_math_h_l150_c3_6613_iffalse := VAR_in24;
     VAR_layer0_node12_MUX_bit_math_h_l150_c3_6613_iftrue := VAR_in25;
     VAR_layer0_node13_MUX_bit_math_h_l161_c3_fd42_iffalse := VAR_in26;
     VAR_layer0_node13_MUX_bit_math_h_l161_c3_fd42_iftrue := VAR_in27;
     VAR_layer0_node14_MUX_bit_math_h_l172_c3_154a_iffalse := VAR_in28;
     VAR_layer0_node14_MUX_bit_math_h_l172_c3_154a_iftrue := VAR_in29;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_0e94_iftrue := VAR_in3;
     VAR_layer0_node15_MUX_bit_math_h_l183_c3_5274_iffalse := VAR_in30;
     VAR_layer0_node15_MUX_bit_math_h_l183_c3_5274_iftrue := VAR_in31;
     VAR_layer0_node16_MUX_bit_math_h_l194_c3_7a7d_iffalse := VAR_in32;
     VAR_layer0_node16_MUX_bit_math_h_l194_c3_7a7d_iftrue := VAR_in33;
     VAR_layer0_node17_MUX_bit_math_h_l205_c3_42ac_iffalse := VAR_in34;
     VAR_layer0_node17_MUX_bit_math_h_l205_c3_42ac_iftrue := VAR_in35;
     VAR_layer0_node18_MUX_bit_math_h_l216_c3_b8f1_iffalse := VAR_in36;
     VAR_layer0_node18_MUX_bit_math_h_l216_c3_b8f1_iftrue := VAR_in37;
     VAR_layer0_node19_MUX_bit_math_h_l227_c3_0b12_iffalse := VAR_in38;
     VAR_layer0_node19_MUX_bit_math_h_l227_c3_0b12_iftrue := VAR_in39;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_e2d9_iffalse := VAR_in4;
     VAR_layer0_node20_MUX_bit_math_h_l238_c3_091e_iffalse := VAR_in40;
     VAR_layer0_node20_MUX_bit_math_h_l238_c3_091e_iftrue := VAR_in41;
     VAR_layer0_node21_MUX_bit_math_h_l249_c3_44d2_iffalse := VAR_in42;
     VAR_layer0_node21_MUX_bit_math_h_l249_c3_44d2_iftrue := VAR_in43;
     VAR_layer0_node22_MUX_bit_math_h_l260_c3_db28_iffalse := VAR_in44;
     VAR_layer0_node22_MUX_bit_math_h_l260_c3_db28_iftrue := VAR_in45;
     VAR_layer0_node23_MUX_bit_math_h_l271_c3_0038_iffalse := VAR_in46;
     VAR_layer0_node23_MUX_bit_math_h_l271_c3_0038_iftrue := VAR_in47;
     VAR_layer0_node24_MUX_bit_math_h_l282_c3_1d56_iffalse := VAR_in48;
     VAR_layer0_node24_MUX_bit_math_h_l282_c3_1d56_iftrue := VAR_in49;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_e2d9_iftrue := VAR_in5;
     VAR_layer0_node25_MUX_bit_math_h_l293_c3_fa3c_iffalse := VAR_in50;
     VAR_layer0_node25_MUX_bit_math_h_l293_c3_fa3c_iftrue := VAR_in51;
     VAR_layer0_node26_MUX_bit_math_h_l304_c3_220e_iffalse := VAR_in52;
     VAR_layer0_node26_MUX_bit_math_h_l304_c3_220e_iftrue := VAR_in53;
     VAR_layer0_node27_MUX_bit_math_h_l315_c3_37d2_iffalse := VAR_in54;
     VAR_layer0_node27_MUX_bit_math_h_l315_c3_37d2_iftrue := VAR_in55;
     VAR_layer0_node28_MUX_bit_math_h_l326_c3_af14_iffalse := VAR_in56;
     VAR_layer0_node28_MUX_bit_math_h_l326_c3_af14_iftrue := VAR_in57;
     VAR_layer0_node29_MUX_bit_math_h_l337_c3_d491_iffalse := VAR_in58;
     VAR_layer0_node29_MUX_bit_math_h_l337_c3_d491_iftrue := VAR_in59;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_edc9_iffalse := VAR_in6;
     VAR_layer0_node30_MUX_bit_math_h_l348_c3_46cf_iffalse := VAR_in60;
     VAR_layer0_node30_MUX_bit_math_h_l348_c3_46cf_iftrue := VAR_in61;
     VAR_layer0_node31_MUX_bit_math_h_l359_c3_1ee6_iffalse := VAR_in62;
     VAR_layer0_node31_MUX_bit_math_h_l359_c3_1ee6_iftrue := VAR_in63;
     VAR_layer0_node32_MUX_bit_math_h_l370_c3_ee39_iffalse := VAR_in64;
     VAR_layer0_node32_MUX_bit_math_h_l370_c3_ee39_iftrue := VAR_in65;
     VAR_layer0_node33_MUX_bit_math_h_l381_c3_f57d_iffalse := VAR_in66;
     VAR_layer0_node33_MUX_bit_math_h_l381_c3_f57d_iftrue := VAR_in67;
     VAR_layer0_node34_MUX_bit_math_h_l392_c3_8d4e_iffalse := VAR_in68;
     VAR_layer0_node34_MUX_bit_math_h_l392_c3_8d4e_iftrue := VAR_in69;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_edc9_iftrue := VAR_in7;
     VAR_layer0_node35_MUX_bit_math_h_l403_c3_fa1f_iffalse := VAR_in70;
     VAR_layer0_node35_MUX_bit_math_h_l403_c3_fa1f_iftrue := VAR_in71;
     VAR_layer0_node36_MUX_bit_math_h_l414_c3_39b4_iffalse := VAR_in72;
     VAR_layer0_node36_MUX_bit_math_h_l414_c3_39b4_iftrue := VAR_in73;
     VAR_layer0_node37_MUX_bit_math_h_l425_c3_3900_iffalse := VAR_in74;
     VAR_layer0_node37_MUX_bit_math_h_l425_c3_3900_iftrue := VAR_in75;
     VAR_layer0_node38_MUX_bit_math_h_l436_c3_bea2_iffalse := VAR_in76;
     VAR_layer0_node38_MUX_bit_math_h_l436_c3_bea2_iftrue := VAR_in77;
     VAR_layer0_node39_MUX_bit_math_h_l447_c3_3acc_iffalse := VAR_in78;
     VAR_layer0_node39_MUX_bit_math_h_l447_c3_3acc_iftrue := VAR_in79;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_f389_iffalse := VAR_in8;
     VAR_layer0_node40_MUX_bit_math_h_l458_c3_f867_iffalse := VAR_in80;
     VAR_layer0_node40_MUX_bit_math_h_l458_c3_f867_iftrue := VAR_in81;
     VAR_layer0_node41_MUX_bit_math_h_l469_c3_2ffe_iffalse := VAR_in82;
     VAR_layer0_node41_MUX_bit_math_h_l469_c3_2ffe_iftrue := VAR_in83;
     VAR_layer0_node42_MUX_bit_math_h_l480_c3_1c62_iffalse := VAR_in84;
     VAR_layer0_node42_MUX_bit_math_h_l480_c3_1c62_iftrue := VAR_in85;
     VAR_layer0_node43_MUX_bit_math_h_l491_c3_7943_iffalse := VAR_in86;
     VAR_layer0_node43_MUX_bit_math_h_l491_c3_7943_iftrue := VAR_in87;
     VAR_layer0_node44_MUX_bit_math_h_l502_c3_15dc_iffalse := VAR_in88;
     VAR_layer0_node44_MUX_bit_math_h_l502_c3_15dc_iftrue := VAR_in89;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_f389_iftrue := VAR_in9;
     VAR_layer0_node45_MUX_bit_math_h_l513_c3_d638_iffalse := VAR_in90;
     VAR_layer0_node45_MUX_bit_math_h_l513_c3_d638_iftrue := VAR_in91;
     VAR_layer0_node46_MUX_bit_math_h_l524_c3_fdc0_iffalse := VAR_in92;
     VAR_layer0_node46_MUX_bit_math_h_l524_c3_fdc0_iftrue := VAR_in93;
     VAR_layer0_node47_MUX_bit_math_h_l535_c3_1640_iffalse := VAR_in94;
     VAR_layer0_node47_MUX_bit_math_h_l535_c3_1640_iftrue := VAR_in95;
     VAR_layer0_node48_MUX_bit_math_h_l546_c3_b0f6_iffalse := VAR_in96;
     VAR_layer0_node48_MUX_bit_math_h_l546_c3_b0f6_iftrue := VAR_in97;
     VAR_layer0_node49_MUX_bit_math_h_l557_c3_adcc_iffalse := VAR_in98;
     VAR_layer0_node49_MUX_bit_math_h_l557_c3_adcc_iftrue := VAR_in99;
     -- uint7_0_0[bit_math_h_l14_c10_5ba9] LATENCY=0
     VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output := uint7_0_0(
     VAR_sel);

     -- uint7_1_1[bit_math_h_l724_c10_ac1d] LATENCY=0
     VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output := uint7_1_1(
     VAR_sel);

     -- uint7_6_6[bit_math_h_l1436_c10_2ac3] LATENCY=0
     VAR_uint7_6_6_bit_math_h_l1436_c10_2ac3_return_output := uint7_6_6(
     VAR_sel);

     -- uint7_2_2[bit_math_h_l1082_c10_87dc] LATENCY=0
     VAR_uint7_2_2_bit_math_h_l1082_c10_87dc_return_output := uint7_2_2(
     VAR_sel);

     -- uint7_3_3[bit_math_h_l1264_c10_51ff] LATENCY=0
     VAR_uint7_3_3_bit_math_h_l1264_c10_51ff_return_output := uint7_3_3(
     VAR_sel);

     -- uint7_4_4[bit_math_h_l1358_c10_29af] LATENCY=0
     VAR_uint7_4_4_bit_math_h_l1358_c10_29af_return_output := uint7_4_4(
     VAR_sel);

     -- uint7_5_5[bit_math_h_l1408_c10_a313] LATENCY=0
     VAR_uint7_5_5_bit_math_h_l1408_c10_a313_return_output := uint7_5_5(
     VAR_sel);

     -- Submodule level 1
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_ce9b_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node10_MUX_bit_math_h_l128_c3_06f3_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node11_MUX_bit_math_h_l139_c3_dbfc_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node12_MUX_bit_math_h_l150_c3_6613_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node13_MUX_bit_math_h_l161_c3_fd42_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node14_MUX_bit_math_h_l172_c3_154a_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node15_MUX_bit_math_h_l183_c3_5274_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node16_MUX_bit_math_h_l194_c3_7a7d_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node17_MUX_bit_math_h_l205_c3_42ac_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node18_MUX_bit_math_h_l216_c3_b8f1_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node19_MUX_bit_math_h_l227_c3_0b12_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_0e94_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node20_MUX_bit_math_h_l238_c3_091e_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node21_MUX_bit_math_h_l249_c3_44d2_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node22_MUX_bit_math_h_l260_c3_db28_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node23_MUX_bit_math_h_l271_c3_0038_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node24_MUX_bit_math_h_l282_c3_1d56_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node25_MUX_bit_math_h_l293_c3_fa3c_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node26_MUX_bit_math_h_l304_c3_220e_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node27_MUX_bit_math_h_l315_c3_37d2_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node28_MUX_bit_math_h_l326_c3_af14_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node29_MUX_bit_math_h_l337_c3_d491_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_e2d9_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node30_MUX_bit_math_h_l348_c3_46cf_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node31_MUX_bit_math_h_l359_c3_1ee6_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node32_MUX_bit_math_h_l370_c3_ee39_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node33_MUX_bit_math_h_l381_c3_f57d_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node34_MUX_bit_math_h_l392_c3_8d4e_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node35_MUX_bit_math_h_l403_c3_fa1f_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node36_MUX_bit_math_h_l414_c3_39b4_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node37_MUX_bit_math_h_l425_c3_3900_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node38_MUX_bit_math_h_l436_c3_bea2_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node39_MUX_bit_math_h_l447_c3_3acc_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_edc9_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node40_MUX_bit_math_h_l458_c3_f867_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node41_MUX_bit_math_h_l469_c3_2ffe_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node42_MUX_bit_math_h_l480_c3_1c62_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node43_MUX_bit_math_h_l491_c3_7943_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node44_MUX_bit_math_h_l502_c3_15dc_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node45_MUX_bit_math_h_l513_c3_d638_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node46_MUX_bit_math_h_l524_c3_fdc0_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node47_MUX_bit_math_h_l535_c3_1640_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node48_MUX_bit_math_h_l546_c3_b0f6_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node49_MUX_bit_math_h_l557_c3_adcc_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_f389_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node50_MUX_bit_math_h_l568_c3_e90e_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node51_MUX_bit_math_h_l579_c3_221f_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node52_MUX_bit_math_h_l590_c3_70e0_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node53_MUX_bit_math_h_l601_c3_e235_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node54_MUX_bit_math_h_l612_c3_f982_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node55_MUX_bit_math_h_l623_c3_bc3d_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node56_MUX_bit_math_h_l634_c3_8e72_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node57_MUX_bit_math_h_l645_c3_0789_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node58_MUX_bit_math_h_l656_c3_d346_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node59_MUX_bit_math_h_l667_c3_d31e_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_d655_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node60_MUX_bit_math_h_l678_c3_e120_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node61_MUX_bit_math_h_l689_c3_a1a2_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node62_MUX_bit_math_h_l700_c3_4595_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node63_MUX_bit_math_h_l711_c3_c6ab_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_5cd3_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_5030_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node8_MUX_bit_math_h_l106_c3_32cb_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer0_node9_MUX_bit_math_h_l117_c3_4b42_cond := VAR_uint7_0_0_bit_math_h_l14_c10_5ba9_return_output;
     VAR_layer1_node0_MUX_bit_math_h_l728_c3_4268_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node10_MUX_bit_math_h_l838_c3_8a99_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node11_MUX_bit_math_h_l849_c3_e0a5_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node12_MUX_bit_math_h_l860_c3_53b9_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node13_MUX_bit_math_h_l871_c3_672a_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node14_MUX_bit_math_h_l882_c3_2725_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node15_MUX_bit_math_h_l893_c3_b457_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node16_MUX_bit_math_h_l904_c3_8832_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node17_MUX_bit_math_h_l915_c3_0128_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node18_MUX_bit_math_h_l926_c3_a8cf_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node19_MUX_bit_math_h_l937_c3_3d6b_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l739_c3_ff28_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node20_MUX_bit_math_h_l948_c3_331f_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node21_MUX_bit_math_h_l959_c3_32d5_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node22_MUX_bit_math_h_l970_c3_56f9_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node23_MUX_bit_math_h_l981_c3_251b_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node24_MUX_bit_math_h_l992_c3_a508_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node28_MUX_bit_math_h_l1036_c3_064f_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node29_MUX_bit_math_h_l1047_c3_e950_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l750_c3_543f_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node30_MUX_bit_math_h_l1058_c3_fdae_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node31_MUX_bit_math_h_l1069_c3_6030_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l761_c3_5c18_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node4_MUX_bit_math_h_l772_c3_a66b_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node5_MUX_bit_math_h_l783_c3_6db3_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node6_MUX_bit_math_h_l794_c3_4c59_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node7_MUX_bit_math_h_l805_c3_502f_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node8_MUX_bit_math_h_l816_c3_1eec_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer1_node9_MUX_bit_math_h_l827_c3_d105_cond := VAR_uint7_1_1_bit_math_h_l724_c10_ac1d_return_output;
     VAR_layer2_node0_MUX_bit_math_h_l1086_c3_122d_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_87dc_return_output;
     VAR_layer2_node10_MUX_bit_math_h_l1196_c3_1666_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_87dc_return_output;
     VAR_layer2_node11_MUX_bit_math_h_l1207_c3_b8de_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_87dc_return_output;
     VAR_layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_87dc_return_output;
     VAR_layer2_node13_MUX_bit_math_h_l1229_c3_d585_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_87dc_return_output;
     VAR_layer2_node14_MUX_bit_math_h_l1240_c3_beb5_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_87dc_return_output;
     VAR_layer2_node15_MUX_bit_math_h_l1251_c3_7550_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_87dc_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_87dc_return_output;
     VAR_layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_87dc_return_output;
     VAR_layer2_node3_MUX_bit_math_h_l1119_c3_946d_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_87dc_return_output;
     VAR_layer2_node4_MUX_bit_math_h_l1130_c3_1f93_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_87dc_return_output;
     VAR_layer2_node5_MUX_bit_math_h_l1141_c3_1425_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_87dc_return_output;
     VAR_layer2_node6_MUX_bit_math_h_l1152_c3_008a_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_87dc_return_output;
     VAR_layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_87dc_return_output;
     VAR_layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_87dc_return_output;
     VAR_layer2_node9_MUX_bit_math_h_l1185_c3_98c3_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_87dc_return_output;
     VAR_layer3_node0_MUX_bit_math_h_l1268_c3_302d_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_51ff_return_output;
     VAR_layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_51ff_return_output;
     VAR_layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_51ff_return_output;
     VAR_layer3_node3_MUX_bit_math_h_l1301_c3_84c3_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_51ff_return_output;
     VAR_layer3_node4_MUX_bit_math_h_l1312_c3_8c96_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_51ff_return_output;
     VAR_layer3_node5_MUX_bit_math_h_l1323_c3_57ee_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_51ff_return_output;
     VAR_layer3_node6_MUX_bit_math_h_l1334_c3_f24c_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_51ff_return_output;
     VAR_layer3_node7_MUX_bit_math_h_l1345_c3_c68c_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_51ff_return_output;
     VAR_layer4_node0_MUX_bit_math_h_l1362_c3_a122_cond := VAR_uint7_4_4_bit_math_h_l1358_c10_29af_return_output;
     VAR_layer4_node1_MUX_bit_math_h_l1373_c3_c86f_cond := VAR_uint7_4_4_bit_math_h_l1358_c10_29af_return_output;
     VAR_layer4_node2_MUX_bit_math_h_l1384_c3_76f0_cond := VAR_uint7_4_4_bit_math_h_l1358_c10_29af_return_output;
     VAR_layer4_node3_MUX_bit_math_h_l1395_c3_5649_cond := VAR_uint7_4_4_bit_math_h_l1358_c10_29af_return_output;
     VAR_layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_cond := VAR_uint7_5_5_bit_math_h_l1408_c10_a313_return_output;
     VAR_layer5_node1_MUX_bit_math_h_l1423_c3_d92a_cond := VAR_uint7_5_5_bit_math_h_l1408_c10_a313_return_output;
     VAR_layer6_node0_MUX_bit_math_h_l1440_c3_43c9_cond := VAR_uint7_6_6_bit_math_h_l1436_c10_2ac3_return_output;
     -- layer0_node45_MUX[bit_math_h_l513_c3_d638] LATENCY=0
     -- Inputs
     layer0_node45_MUX_bit_math_h_l513_c3_d638_cond <= VAR_layer0_node45_MUX_bit_math_h_l513_c3_d638_cond;
     layer0_node45_MUX_bit_math_h_l513_c3_d638_iftrue <= VAR_layer0_node45_MUX_bit_math_h_l513_c3_d638_iftrue;
     layer0_node45_MUX_bit_math_h_l513_c3_d638_iffalse <= VAR_layer0_node45_MUX_bit_math_h_l513_c3_d638_iffalse;
     -- Outputs
     VAR_layer0_node45_MUX_bit_math_h_l513_c3_d638_return_output := layer0_node45_MUX_bit_math_h_l513_c3_d638_return_output;

     -- layer0_node11_MUX[bit_math_h_l139_c3_dbfc] LATENCY=0
     -- Inputs
     layer0_node11_MUX_bit_math_h_l139_c3_dbfc_cond <= VAR_layer0_node11_MUX_bit_math_h_l139_c3_dbfc_cond;
     layer0_node11_MUX_bit_math_h_l139_c3_dbfc_iftrue <= VAR_layer0_node11_MUX_bit_math_h_l139_c3_dbfc_iftrue;
     layer0_node11_MUX_bit_math_h_l139_c3_dbfc_iffalse <= VAR_layer0_node11_MUX_bit_math_h_l139_c3_dbfc_iffalse;
     -- Outputs
     VAR_layer0_node11_MUX_bit_math_h_l139_c3_dbfc_return_output := layer0_node11_MUX_bit_math_h_l139_c3_dbfc_return_output;

     -- layer0_node58_MUX[bit_math_h_l656_c3_d346] LATENCY=0
     -- Inputs
     layer0_node58_MUX_bit_math_h_l656_c3_d346_cond <= VAR_layer0_node58_MUX_bit_math_h_l656_c3_d346_cond;
     layer0_node58_MUX_bit_math_h_l656_c3_d346_iftrue <= VAR_layer0_node58_MUX_bit_math_h_l656_c3_d346_iftrue;
     layer0_node58_MUX_bit_math_h_l656_c3_d346_iffalse <= VAR_layer0_node58_MUX_bit_math_h_l656_c3_d346_iffalse;
     -- Outputs
     VAR_layer0_node58_MUX_bit_math_h_l656_c3_d346_return_output := layer0_node58_MUX_bit_math_h_l656_c3_d346_return_output;

     -- layer0_node9_MUX[bit_math_h_l117_c3_4b42] LATENCY=0
     -- Inputs
     layer0_node9_MUX_bit_math_h_l117_c3_4b42_cond <= VAR_layer0_node9_MUX_bit_math_h_l117_c3_4b42_cond;
     layer0_node9_MUX_bit_math_h_l117_c3_4b42_iftrue <= VAR_layer0_node9_MUX_bit_math_h_l117_c3_4b42_iftrue;
     layer0_node9_MUX_bit_math_h_l117_c3_4b42_iffalse <= VAR_layer0_node9_MUX_bit_math_h_l117_c3_4b42_iffalse;
     -- Outputs
     VAR_layer0_node9_MUX_bit_math_h_l117_c3_4b42_return_output := layer0_node9_MUX_bit_math_h_l117_c3_4b42_return_output;

     -- layer0_node12_MUX[bit_math_h_l150_c3_6613] LATENCY=0
     -- Inputs
     layer0_node12_MUX_bit_math_h_l150_c3_6613_cond <= VAR_layer0_node12_MUX_bit_math_h_l150_c3_6613_cond;
     layer0_node12_MUX_bit_math_h_l150_c3_6613_iftrue <= VAR_layer0_node12_MUX_bit_math_h_l150_c3_6613_iftrue;
     layer0_node12_MUX_bit_math_h_l150_c3_6613_iffalse <= VAR_layer0_node12_MUX_bit_math_h_l150_c3_6613_iffalse;
     -- Outputs
     VAR_layer0_node12_MUX_bit_math_h_l150_c3_6613_return_output := layer0_node12_MUX_bit_math_h_l150_c3_6613_return_output;

     -- layer0_node27_MUX[bit_math_h_l315_c3_37d2] LATENCY=0
     -- Inputs
     layer0_node27_MUX_bit_math_h_l315_c3_37d2_cond <= VAR_layer0_node27_MUX_bit_math_h_l315_c3_37d2_cond;
     layer0_node27_MUX_bit_math_h_l315_c3_37d2_iftrue <= VAR_layer0_node27_MUX_bit_math_h_l315_c3_37d2_iftrue;
     layer0_node27_MUX_bit_math_h_l315_c3_37d2_iffalse <= VAR_layer0_node27_MUX_bit_math_h_l315_c3_37d2_iffalse;
     -- Outputs
     VAR_layer0_node27_MUX_bit_math_h_l315_c3_37d2_return_output := layer0_node27_MUX_bit_math_h_l315_c3_37d2_return_output;

     -- layer0_node61_MUX[bit_math_h_l689_c3_a1a2] LATENCY=0
     -- Inputs
     layer0_node61_MUX_bit_math_h_l689_c3_a1a2_cond <= VAR_layer0_node61_MUX_bit_math_h_l689_c3_a1a2_cond;
     layer0_node61_MUX_bit_math_h_l689_c3_a1a2_iftrue <= VAR_layer0_node61_MUX_bit_math_h_l689_c3_a1a2_iftrue;
     layer0_node61_MUX_bit_math_h_l689_c3_a1a2_iffalse <= VAR_layer0_node61_MUX_bit_math_h_l689_c3_a1a2_iffalse;
     -- Outputs
     VAR_layer0_node61_MUX_bit_math_h_l689_c3_a1a2_return_output := layer0_node61_MUX_bit_math_h_l689_c3_a1a2_return_output;

     -- layer0_node5_MUX[bit_math_h_l73_c3_d655] LATENCY=0
     -- Inputs
     layer0_node5_MUX_bit_math_h_l73_c3_d655_cond <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_d655_cond;
     layer0_node5_MUX_bit_math_h_l73_c3_d655_iftrue <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_d655_iftrue;
     layer0_node5_MUX_bit_math_h_l73_c3_d655_iffalse <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_d655_iffalse;
     -- Outputs
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_d655_return_output := layer0_node5_MUX_bit_math_h_l73_c3_d655_return_output;

     -- layer0_node33_MUX[bit_math_h_l381_c3_f57d] LATENCY=0
     -- Inputs
     layer0_node33_MUX_bit_math_h_l381_c3_f57d_cond <= VAR_layer0_node33_MUX_bit_math_h_l381_c3_f57d_cond;
     layer0_node33_MUX_bit_math_h_l381_c3_f57d_iftrue <= VAR_layer0_node33_MUX_bit_math_h_l381_c3_f57d_iftrue;
     layer0_node33_MUX_bit_math_h_l381_c3_f57d_iffalse <= VAR_layer0_node33_MUX_bit_math_h_l381_c3_f57d_iffalse;
     -- Outputs
     VAR_layer0_node33_MUX_bit_math_h_l381_c3_f57d_return_output := layer0_node33_MUX_bit_math_h_l381_c3_f57d_return_output;

     -- layer0_node34_MUX[bit_math_h_l392_c3_8d4e] LATENCY=0
     -- Inputs
     layer0_node34_MUX_bit_math_h_l392_c3_8d4e_cond <= VAR_layer0_node34_MUX_bit_math_h_l392_c3_8d4e_cond;
     layer0_node34_MUX_bit_math_h_l392_c3_8d4e_iftrue <= VAR_layer0_node34_MUX_bit_math_h_l392_c3_8d4e_iftrue;
     layer0_node34_MUX_bit_math_h_l392_c3_8d4e_iffalse <= VAR_layer0_node34_MUX_bit_math_h_l392_c3_8d4e_iffalse;
     -- Outputs
     VAR_layer0_node34_MUX_bit_math_h_l392_c3_8d4e_return_output := layer0_node34_MUX_bit_math_h_l392_c3_8d4e_return_output;

     -- layer0_node43_MUX[bit_math_h_l491_c3_7943] LATENCY=0
     -- Inputs
     layer0_node43_MUX_bit_math_h_l491_c3_7943_cond <= VAR_layer0_node43_MUX_bit_math_h_l491_c3_7943_cond;
     layer0_node43_MUX_bit_math_h_l491_c3_7943_iftrue <= VAR_layer0_node43_MUX_bit_math_h_l491_c3_7943_iftrue;
     layer0_node43_MUX_bit_math_h_l491_c3_7943_iffalse <= VAR_layer0_node43_MUX_bit_math_h_l491_c3_7943_iffalse;
     -- Outputs
     VAR_layer0_node43_MUX_bit_math_h_l491_c3_7943_return_output := layer0_node43_MUX_bit_math_h_l491_c3_7943_return_output;

     -- layer0_node54_MUX[bit_math_h_l612_c3_f982] LATENCY=0
     -- Inputs
     layer0_node54_MUX_bit_math_h_l612_c3_f982_cond <= VAR_layer0_node54_MUX_bit_math_h_l612_c3_f982_cond;
     layer0_node54_MUX_bit_math_h_l612_c3_f982_iftrue <= VAR_layer0_node54_MUX_bit_math_h_l612_c3_f982_iftrue;
     layer0_node54_MUX_bit_math_h_l612_c3_f982_iffalse <= VAR_layer0_node54_MUX_bit_math_h_l612_c3_f982_iffalse;
     -- Outputs
     VAR_layer0_node54_MUX_bit_math_h_l612_c3_f982_return_output := layer0_node54_MUX_bit_math_h_l612_c3_f982_return_output;

     -- layer0_node59_MUX[bit_math_h_l667_c3_d31e] LATENCY=0
     -- Inputs
     layer0_node59_MUX_bit_math_h_l667_c3_d31e_cond <= VAR_layer0_node59_MUX_bit_math_h_l667_c3_d31e_cond;
     layer0_node59_MUX_bit_math_h_l667_c3_d31e_iftrue <= VAR_layer0_node59_MUX_bit_math_h_l667_c3_d31e_iftrue;
     layer0_node59_MUX_bit_math_h_l667_c3_d31e_iffalse <= VAR_layer0_node59_MUX_bit_math_h_l667_c3_d31e_iffalse;
     -- Outputs
     VAR_layer0_node59_MUX_bit_math_h_l667_c3_d31e_return_output := layer0_node59_MUX_bit_math_h_l667_c3_d31e_return_output;

     -- layer0_node10_MUX[bit_math_h_l128_c3_06f3] LATENCY=0
     -- Inputs
     layer0_node10_MUX_bit_math_h_l128_c3_06f3_cond <= VAR_layer0_node10_MUX_bit_math_h_l128_c3_06f3_cond;
     layer0_node10_MUX_bit_math_h_l128_c3_06f3_iftrue <= VAR_layer0_node10_MUX_bit_math_h_l128_c3_06f3_iftrue;
     layer0_node10_MUX_bit_math_h_l128_c3_06f3_iffalse <= VAR_layer0_node10_MUX_bit_math_h_l128_c3_06f3_iffalse;
     -- Outputs
     VAR_layer0_node10_MUX_bit_math_h_l128_c3_06f3_return_output := layer0_node10_MUX_bit_math_h_l128_c3_06f3_return_output;

     -- layer0_node48_MUX[bit_math_h_l546_c3_b0f6] LATENCY=0
     -- Inputs
     layer0_node48_MUX_bit_math_h_l546_c3_b0f6_cond <= VAR_layer0_node48_MUX_bit_math_h_l546_c3_b0f6_cond;
     layer0_node48_MUX_bit_math_h_l546_c3_b0f6_iftrue <= VAR_layer0_node48_MUX_bit_math_h_l546_c3_b0f6_iftrue;
     layer0_node48_MUX_bit_math_h_l546_c3_b0f6_iffalse <= VAR_layer0_node48_MUX_bit_math_h_l546_c3_b0f6_iffalse;
     -- Outputs
     VAR_layer0_node48_MUX_bit_math_h_l546_c3_b0f6_return_output := layer0_node48_MUX_bit_math_h_l546_c3_b0f6_return_output;

     -- layer0_node8_MUX[bit_math_h_l106_c3_32cb] LATENCY=0
     -- Inputs
     layer0_node8_MUX_bit_math_h_l106_c3_32cb_cond <= VAR_layer0_node8_MUX_bit_math_h_l106_c3_32cb_cond;
     layer0_node8_MUX_bit_math_h_l106_c3_32cb_iftrue <= VAR_layer0_node8_MUX_bit_math_h_l106_c3_32cb_iftrue;
     layer0_node8_MUX_bit_math_h_l106_c3_32cb_iffalse <= VAR_layer0_node8_MUX_bit_math_h_l106_c3_32cb_iffalse;
     -- Outputs
     VAR_layer0_node8_MUX_bit_math_h_l106_c3_32cb_return_output := layer0_node8_MUX_bit_math_h_l106_c3_32cb_return_output;

     -- layer0_node51_MUX[bit_math_h_l579_c3_221f] LATENCY=0
     -- Inputs
     layer0_node51_MUX_bit_math_h_l579_c3_221f_cond <= VAR_layer0_node51_MUX_bit_math_h_l579_c3_221f_cond;
     layer0_node51_MUX_bit_math_h_l579_c3_221f_iftrue <= VAR_layer0_node51_MUX_bit_math_h_l579_c3_221f_iftrue;
     layer0_node51_MUX_bit_math_h_l579_c3_221f_iffalse <= VAR_layer0_node51_MUX_bit_math_h_l579_c3_221f_iffalse;
     -- Outputs
     VAR_layer0_node51_MUX_bit_math_h_l579_c3_221f_return_output := layer0_node51_MUX_bit_math_h_l579_c3_221f_return_output;

     -- layer0_node29_MUX[bit_math_h_l337_c3_d491] LATENCY=0
     -- Inputs
     layer0_node29_MUX_bit_math_h_l337_c3_d491_cond <= VAR_layer0_node29_MUX_bit_math_h_l337_c3_d491_cond;
     layer0_node29_MUX_bit_math_h_l337_c3_d491_iftrue <= VAR_layer0_node29_MUX_bit_math_h_l337_c3_d491_iftrue;
     layer0_node29_MUX_bit_math_h_l337_c3_d491_iffalse <= VAR_layer0_node29_MUX_bit_math_h_l337_c3_d491_iffalse;
     -- Outputs
     VAR_layer0_node29_MUX_bit_math_h_l337_c3_d491_return_output := layer0_node29_MUX_bit_math_h_l337_c3_d491_return_output;

     -- layer0_node25_MUX[bit_math_h_l293_c3_fa3c] LATENCY=0
     -- Inputs
     layer0_node25_MUX_bit_math_h_l293_c3_fa3c_cond <= VAR_layer0_node25_MUX_bit_math_h_l293_c3_fa3c_cond;
     layer0_node25_MUX_bit_math_h_l293_c3_fa3c_iftrue <= VAR_layer0_node25_MUX_bit_math_h_l293_c3_fa3c_iftrue;
     layer0_node25_MUX_bit_math_h_l293_c3_fa3c_iffalse <= VAR_layer0_node25_MUX_bit_math_h_l293_c3_fa3c_iffalse;
     -- Outputs
     VAR_layer0_node25_MUX_bit_math_h_l293_c3_fa3c_return_output := layer0_node25_MUX_bit_math_h_l293_c3_fa3c_return_output;

     -- layer0_node52_MUX[bit_math_h_l590_c3_70e0] LATENCY=0
     -- Inputs
     layer0_node52_MUX_bit_math_h_l590_c3_70e0_cond <= VAR_layer0_node52_MUX_bit_math_h_l590_c3_70e0_cond;
     layer0_node52_MUX_bit_math_h_l590_c3_70e0_iftrue <= VAR_layer0_node52_MUX_bit_math_h_l590_c3_70e0_iftrue;
     layer0_node52_MUX_bit_math_h_l590_c3_70e0_iffalse <= VAR_layer0_node52_MUX_bit_math_h_l590_c3_70e0_iffalse;
     -- Outputs
     VAR_layer0_node52_MUX_bit_math_h_l590_c3_70e0_return_output := layer0_node52_MUX_bit_math_h_l590_c3_70e0_return_output;

     -- layer0_node42_MUX[bit_math_h_l480_c3_1c62] LATENCY=0
     -- Inputs
     layer0_node42_MUX_bit_math_h_l480_c3_1c62_cond <= VAR_layer0_node42_MUX_bit_math_h_l480_c3_1c62_cond;
     layer0_node42_MUX_bit_math_h_l480_c3_1c62_iftrue <= VAR_layer0_node42_MUX_bit_math_h_l480_c3_1c62_iftrue;
     layer0_node42_MUX_bit_math_h_l480_c3_1c62_iffalse <= VAR_layer0_node42_MUX_bit_math_h_l480_c3_1c62_iffalse;
     -- Outputs
     VAR_layer0_node42_MUX_bit_math_h_l480_c3_1c62_return_output := layer0_node42_MUX_bit_math_h_l480_c3_1c62_return_output;

     -- layer0_node17_MUX[bit_math_h_l205_c3_42ac] LATENCY=0
     -- Inputs
     layer0_node17_MUX_bit_math_h_l205_c3_42ac_cond <= VAR_layer0_node17_MUX_bit_math_h_l205_c3_42ac_cond;
     layer0_node17_MUX_bit_math_h_l205_c3_42ac_iftrue <= VAR_layer0_node17_MUX_bit_math_h_l205_c3_42ac_iftrue;
     layer0_node17_MUX_bit_math_h_l205_c3_42ac_iffalse <= VAR_layer0_node17_MUX_bit_math_h_l205_c3_42ac_iffalse;
     -- Outputs
     VAR_layer0_node17_MUX_bit_math_h_l205_c3_42ac_return_output := layer0_node17_MUX_bit_math_h_l205_c3_42ac_return_output;

     -- layer0_node26_MUX[bit_math_h_l304_c3_220e] LATENCY=0
     -- Inputs
     layer0_node26_MUX_bit_math_h_l304_c3_220e_cond <= VAR_layer0_node26_MUX_bit_math_h_l304_c3_220e_cond;
     layer0_node26_MUX_bit_math_h_l304_c3_220e_iftrue <= VAR_layer0_node26_MUX_bit_math_h_l304_c3_220e_iftrue;
     layer0_node26_MUX_bit_math_h_l304_c3_220e_iffalse <= VAR_layer0_node26_MUX_bit_math_h_l304_c3_220e_iffalse;
     -- Outputs
     VAR_layer0_node26_MUX_bit_math_h_l304_c3_220e_return_output := layer0_node26_MUX_bit_math_h_l304_c3_220e_return_output;

     -- layer0_node63_MUX[bit_math_h_l711_c3_c6ab] LATENCY=0
     -- Inputs
     layer0_node63_MUX_bit_math_h_l711_c3_c6ab_cond <= VAR_layer0_node63_MUX_bit_math_h_l711_c3_c6ab_cond;
     layer0_node63_MUX_bit_math_h_l711_c3_c6ab_iftrue <= VAR_layer0_node63_MUX_bit_math_h_l711_c3_c6ab_iftrue;
     layer0_node63_MUX_bit_math_h_l711_c3_c6ab_iffalse <= VAR_layer0_node63_MUX_bit_math_h_l711_c3_c6ab_iffalse;
     -- Outputs
     VAR_layer0_node63_MUX_bit_math_h_l711_c3_c6ab_return_output := layer0_node63_MUX_bit_math_h_l711_c3_c6ab_return_output;

     -- layer0_node31_MUX[bit_math_h_l359_c3_1ee6] LATENCY=0
     -- Inputs
     layer0_node31_MUX_bit_math_h_l359_c3_1ee6_cond <= VAR_layer0_node31_MUX_bit_math_h_l359_c3_1ee6_cond;
     layer0_node31_MUX_bit_math_h_l359_c3_1ee6_iftrue <= VAR_layer0_node31_MUX_bit_math_h_l359_c3_1ee6_iftrue;
     layer0_node31_MUX_bit_math_h_l359_c3_1ee6_iffalse <= VAR_layer0_node31_MUX_bit_math_h_l359_c3_1ee6_iffalse;
     -- Outputs
     VAR_layer0_node31_MUX_bit_math_h_l359_c3_1ee6_return_output := layer0_node31_MUX_bit_math_h_l359_c3_1ee6_return_output;

     -- layer0_node60_MUX[bit_math_h_l678_c3_e120] LATENCY=0
     -- Inputs
     layer0_node60_MUX_bit_math_h_l678_c3_e120_cond <= VAR_layer0_node60_MUX_bit_math_h_l678_c3_e120_cond;
     layer0_node60_MUX_bit_math_h_l678_c3_e120_iftrue <= VAR_layer0_node60_MUX_bit_math_h_l678_c3_e120_iftrue;
     layer0_node60_MUX_bit_math_h_l678_c3_e120_iffalse <= VAR_layer0_node60_MUX_bit_math_h_l678_c3_e120_iffalse;
     -- Outputs
     VAR_layer0_node60_MUX_bit_math_h_l678_c3_e120_return_output := layer0_node60_MUX_bit_math_h_l678_c3_e120_return_output;

     -- layer0_node13_MUX[bit_math_h_l161_c3_fd42] LATENCY=0
     -- Inputs
     layer0_node13_MUX_bit_math_h_l161_c3_fd42_cond <= VAR_layer0_node13_MUX_bit_math_h_l161_c3_fd42_cond;
     layer0_node13_MUX_bit_math_h_l161_c3_fd42_iftrue <= VAR_layer0_node13_MUX_bit_math_h_l161_c3_fd42_iftrue;
     layer0_node13_MUX_bit_math_h_l161_c3_fd42_iffalse <= VAR_layer0_node13_MUX_bit_math_h_l161_c3_fd42_iffalse;
     -- Outputs
     VAR_layer0_node13_MUX_bit_math_h_l161_c3_fd42_return_output := layer0_node13_MUX_bit_math_h_l161_c3_fd42_return_output;

     -- layer0_node53_MUX[bit_math_h_l601_c3_e235] LATENCY=0
     -- Inputs
     layer0_node53_MUX_bit_math_h_l601_c3_e235_cond <= VAR_layer0_node53_MUX_bit_math_h_l601_c3_e235_cond;
     layer0_node53_MUX_bit_math_h_l601_c3_e235_iftrue <= VAR_layer0_node53_MUX_bit_math_h_l601_c3_e235_iftrue;
     layer0_node53_MUX_bit_math_h_l601_c3_e235_iffalse <= VAR_layer0_node53_MUX_bit_math_h_l601_c3_e235_iffalse;
     -- Outputs
     VAR_layer0_node53_MUX_bit_math_h_l601_c3_e235_return_output := layer0_node53_MUX_bit_math_h_l601_c3_e235_return_output;

     -- layer0_node28_MUX[bit_math_h_l326_c3_af14] LATENCY=0
     -- Inputs
     layer0_node28_MUX_bit_math_h_l326_c3_af14_cond <= VAR_layer0_node28_MUX_bit_math_h_l326_c3_af14_cond;
     layer0_node28_MUX_bit_math_h_l326_c3_af14_iftrue <= VAR_layer0_node28_MUX_bit_math_h_l326_c3_af14_iftrue;
     layer0_node28_MUX_bit_math_h_l326_c3_af14_iffalse <= VAR_layer0_node28_MUX_bit_math_h_l326_c3_af14_iffalse;
     -- Outputs
     VAR_layer0_node28_MUX_bit_math_h_l326_c3_af14_return_output := layer0_node28_MUX_bit_math_h_l326_c3_af14_return_output;

     -- layer0_node55_MUX[bit_math_h_l623_c3_bc3d] LATENCY=0
     -- Inputs
     layer0_node55_MUX_bit_math_h_l623_c3_bc3d_cond <= VAR_layer0_node55_MUX_bit_math_h_l623_c3_bc3d_cond;
     layer0_node55_MUX_bit_math_h_l623_c3_bc3d_iftrue <= VAR_layer0_node55_MUX_bit_math_h_l623_c3_bc3d_iftrue;
     layer0_node55_MUX_bit_math_h_l623_c3_bc3d_iffalse <= VAR_layer0_node55_MUX_bit_math_h_l623_c3_bc3d_iffalse;
     -- Outputs
     VAR_layer0_node55_MUX_bit_math_h_l623_c3_bc3d_return_output := layer0_node55_MUX_bit_math_h_l623_c3_bc3d_return_output;

     -- layer0_node19_MUX[bit_math_h_l227_c3_0b12] LATENCY=0
     -- Inputs
     layer0_node19_MUX_bit_math_h_l227_c3_0b12_cond <= VAR_layer0_node19_MUX_bit_math_h_l227_c3_0b12_cond;
     layer0_node19_MUX_bit_math_h_l227_c3_0b12_iftrue <= VAR_layer0_node19_MUX_bit_math_h_l227_c3_0b12_iftrue;
     layer0_node19_MUX_bit_math_h_l227_c3_0b12_iffalse <= VAR_layer0_node19_MUX_bit_math_h_l227_c3_0b12_iffalse;
     -- Outputs
     VAR_layer0_node19_MUX_bit_math_h_l227_c3_0b12_return_output := layer0_node19_MUX_bit_math_h_l227_c3_0b12_return_output;

     -- layer0_node50_MUX[bit_math_h_l568_c3_e90e] LATENCY=0
     -- Inputs
     layer0_node50_MUX_bit_math_h_l568_c3_e90e_cond <= VAR_layer0_node50_MUX_bit_math_h_l568_c3_e90e_cond;
     layer0_node50_MUX_bit_math_h_l568_c3_e90e_iftrue <= VAR_layer0_node50_MUX_bit_math_h_l568_c3_e90e_iftrue;
     layer0_node50_MUX_bit_math_h_l568_c3_e90e_iffalse <= VAR_layer0_node50_MUX_bit_math_h_l568_c3_e90e_iffalse;
     -- Outputs
     VAR_layer0_node50_MUX_bit_math_h_l568_c3_e90e_return_output := layer0_node50_MUX_bit_math_h_l568_c3_e90e_return_output;

     -- layer0_node46_MUX[bit_math_h_l524_c3_fdc0] LATENCY=0
     -- Inputs
     layer0_node46_MUX_bit_math_h_l524_c3_fdc0_cond <= VAR_layer0_node46_MUX_bit_math_h_l524_c3_fdc0_cond;
     layer0_node46_MUX_bit_math_h_l524_c3_fdc0_iftrue <= VAR_layer0_node46_MUX_bit_math_h_l524_c3_fdc0_iftrue;
     layer0_node46_MUX_bit_math_h_l524_c3_fdc0_iffalse <= VAR_layer0_node46_MUX_bit_math_h_l524_c3_fdc0_iffalse;
     -- Outputs
     VAR_layer0_node46_MUX_bit_math_h_l524_c3_fdc0_return_output := layer0_node46_MUX_bit_math_h_l524_c3_fdc0_return_output;

     -- layer0_node4_MUX[bit_math_h_l62_c3_f389] LATENCY=0
     -- Inputs
     layer0_node4_MUX_bit_math_h_l62_c3_f389_cond <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_f389_cond;
     layer0_node4_MUX_bit_math_h_l62_c3_f389_iftrue <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_f389_iftrue;
     layer0_node4_MUX_bit_math_h_l62_c3_f389_iffalse <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_f389_iffalse;
     -- Outputs
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_f389_return_output := layer0_node4_MUX_bit_math_h_l62_c3_f389_return_output;

     -- layer0_node47_MUX[bit_math_h_l535_c3_1640] LATENCY=0
     -- Inputs
     layer0_node47_MUX_bit_math_h_l535_c3_1640_cond <= VAR_layer0_node47_MUX_bit_math_h_l535_c3_1640_cond;
     layer0_node47_MUX_bit_math_h_l535_c3_1640_iftrue <= VAR_layer0_node47_MUX_bit_math_h_l535_c3_1640_iftrue;
     layer0_node47_MUX_bit_math_h_l535_c3_1640_iffalse <= VAR_layer0_node47_MUX_bit_math_h_l535_c3_1640_iffalse;
     -- Outputs
     VAR_layer0_node47_MUX_bit_math_h_l535_c3_1640_return_output := layer0_node47_MUX_bit_math_h_l535_c3_1640_return_output;

     -- layer0_node57_MUX[bit_math_h_l645_c3_0789] LATENCY=0
     -- Inputs
     layer0_node57_MUX_bit_math_h_l645_c3_0789_cond <= VAR_layer0_node57_MUX_bit_math_h_l645_c3_0789_cond;
     layer0_node57_MUX_bit_math_h_l645_c3_0789_iftrue <= VAR_layer0_node57_MUX_bit_math_h_l645_c3_0789_iftrue;
     layer0_node57_MUX_bit_math_h_l645_c3_0789_iffalse <= VAR_layer0_node57_MUX_bit_math_h_l645_c3_0789_iffalse;
     -- Outputs
     VAR_layer0_node57_MUX_bit_math_h_l645_c3_0789_return_output := layer0_node57_MUX_bit_math_h_l645_c3_0789_return_output;

     -- layer0_node21_MUX[bit_math_h_l249_c3_44d2] LATENCY=0
     -- Inputs
     layer0_node21_MUX_bit_math_h_l249_c3_44d2_cond <= VAR_layer0_node21_MUX_bit_math_h_l249_c3_44d2_cond;
     layer0_node21_MUX_bit_math_h_l249_c3_44d2_iftrue <= VAR_layer0_node21_MUX_bit_math_h_l249_c3_44d2_iftrue;
     layer0_node21_MUX_bit_math_h_l249_c3_44d2_iffalse <= VAR_layer0_node21_MUX_bit_math_h_l249_c3_44d2_iffalse;
     -- Outputs
     VAR_layer0_node21_MUX_bit_math_h_l249_c3_44d2_return_output := layer0_node21_MUX_bit_math_h_l249_c3_44d2_return_output;

     -- layer0_node32_MUX[bit_math_h_l370_c3_ee39] LATENCY=0
     -- Inputs
     layer0_node32_MUX_bit_math_h_l370_c3_ee39_cond <= VAR_layer0_node32_MUX_bit_math_h_l370_c3_ee39_cond;
     layer0_node32_MUX_bit_math_h_l370_c3_ee39_iftrue <= VAR_layer0_node32_MUX_bit_math_h_l370_c3_ee39_iftrue;
     layer0_node32_MUX_bit_math_h_l370_c3_ee39_iffalse <= VAR_layer0_node32_MUX_bit_math_h_l370_c3_ee39_iffalse;
     -- Outputs
     VAR_layer0_node32_MUX_bit_math_h_l370_c3_ee39_return_output := layer0_node32_MUX_bit_math_h_l370_c3_ee39_return_output;

     -- layer0_node2_MUX[bit_math_h_l40_c3_e2d9] LATENCY=0
     -- Inputs
     layer0_node2_MUX_bit_math_h_l40_c3_e2d9_cond <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_e2d9_cond;
     layer0_node2_MUX_bit_math_h_l40_c3_e2d9_iftrue <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_e2d9_iftrue;
     layer0_node2_MUX_bit_math_h_l40_c3_e2d9_iffalse <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_e2d9_iffalse;
     -- Outputs
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_e2d9_return_output := layer0_node2_MUX_bit_math_h_l40_c3_e2d9_return_output;

     -- layer0_node35_MUX[bit_math_h_l403_c3_fa1f] LATENCY=0
     -- Inputs
     layer0_node35_MUX_bit_math_h_l403_c3_fa1f_cond <= VAR_layer0_node35_MUX_bit_math_h_l403_c3_fa1f_cond;
     layer0_node35_MUX_bit_math_h_l403_c3_fa1f_iftrue <= VAR_layer0_node35_MUX_bit_math_h_l403_c3_fa1f_iftrue;
     layer0_node35_MUX_bit_math_h_l403_c3_fa1f_iffalse <= VAR_layer0_node35_MUX_bit_math_h_l403_c3_fa1f_iffalse;
     -- Outputs
     VAR_layer0_node35_MUX_bit_math_h_l403_c3_fa1f_return_output := layer0_node35_MUX_bit_math_h_l403_c3_fa1f_return_output;

     -- layer0_node7_MUX[bit_math_h_l95_c3_5030] LATENCY=0
     -- Inputs
     layer0_node7_MUX_bit_math_h_l95_c3_5030_cond <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_5030_cond;
     layer0_node7_MUX_bit_math_h_l95_c3_5030_iftrue <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_5030_iftrue;
     layer0_node7_MUX_bit_math_h_l95_c3_5030_iffalse <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_5030_iffalse;
     -- Outputs
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_5030_return_output := layer0_node7_MUX_bit_math_h_l95_c3_5030_return_output;

     -- layer0_node6_MUX[bit_math_h_l84_c3_5cd3] LATENCY=0
     -- Inputs
     layer0_node6_MUX_bit_math_h_l84_c3_5cd3_cond <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_5cd3_cond;
     layer0_node6_MUX_bit_math_h_l84_c3_5cd3_iftrue <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_5cd3_iftrue;
     layer0_node6_MUX_bit_math_h_l84_c3_5cd3_iffalse <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_5cd3_iffalse;
     -- Outputs
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_5cd3_return_output := layer0_node6_MUX_bit_math_h_l84_c3_5cd3_return_output;

     -- layer0_node62_MUX[bit_math_h_l700_c3_4595] LATENCY=0
     -- Inputs
     layer0_node62_MUX_bit_math_h_l700_c3_4595_cond <= VAR_layer0_node62_MUX_bit_math_h_l700_c3_4595_cond;
     layer0_node62_MUX_bit_math_h_l700_c3_4595_iftrue <= VAR_layer0_node62_MUX_bit_math_h_l700_c3_4595_iftrue;
     layer0_node62_MUX_bit_math_h_l700_c3_4595_iffalse <= VAR_layer0_node62_MUX_bit_math_h_l700_c3_4595_iffalse;
     -- Outputs
     VAR_layer0_node62_MUX_bit_math_h_l700_c3_4595_return_output := layer0_node62_MUX_bit_math_h_l700_c3_4595_return_output;

     -- layer0_node49_MUX[bit_math_h_l557_c3_adcc] LATENCY=0
     -- Inputs
     layer0_node49_MUX_bit_math_h_l557_c3_adcc_cond <= VAR_layer0_node49_MUX_bit_math_h_l557_c3_adcc_cond;
     layer0_node49_MUX_bit_math_h_l557_c3_adcc_iftrue <= VAR_layer0_node49_MUX_bit_math_h_l557_c3_adcc_iftrue;
     layer0_node49_MUX_bit_math_h_l557_c3_adcc_iffalse <= VAR_layer0_node49_MUX_bit_math_h_l557_c3_adcc_iffalse;
     -- Outputs
     VAR_layer0_node49_MUX_bit_math_h_l557_c3_adcc_return_output := layer0_node49_MUX_bit_math_h_l557_c3_adcc_return_output;

     -- layer0_node36_MUX[bit_math_h_l414_c3_39b4] LATENCY=0
     -- Inputs
     layer0_node36_MUX_bit_math_h_l414_c3_39b4_cond <= VAR_layer0_node36_MUX_bit_math_h_l414_c3_39b4_cond;
     layer0_node36_MUX_bit_math_h_l414_c3_39b4_iftrue <= VAR_layer0_node36_MUX_bit_math_h_l414_c3_39b4_iftrue;
     layer0_node36_MUX_bit_math_h_l414_c3_39b4_iffalse <= VAR_layer0_node36_MUX_bit_math_h_l414_c3_39b4_iffalse;
     -- Outputs
     VAR_layer0_node36_MUX_bit_math_h_l414_c3_39b4_return_output := layer0_node36_MUX_bit_math_h_l414_c3_39b4_return_output;

     -- layer0_node14_MUX[bit_math_h_l172_c3_154a] LATENCY=0
     -- Inputs
     layer0_node14_MUX_bit_math_h_l172_c3_154a_cond <= VAR_layer0_node14_MUX_bit_math_h_l172_c3_154a_cond;
     layer0_node14_MUX_bit_math_h_l172_c3_154a_iftrue <= VAR_layer0_node14_MUX_bit_math_h_l172_c3_154a_iftrue;
     layer0_node14_MUX_bit_math_h_l172_c3_154a_iffalse <= VAR_layer0_node14_MUX_bit_math_h_l172_c3_154a_iffalse;
     -- Outputs
     VAR_layer0_node14_MUX_bit_math_h_l172_c3_154a_return_output := layer0_node14_MUX_bit_math_h_l172_c3_154a_return_output;

     -- layer0_node3_MUX[bit_math_h_l51_c3_edc9] LATENCY=0
     -- Inputs
     layer0_node3_MUX_bit_math_h_l51_c3_edc9_cond <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_edc9_cond;
     layer0_node3_MUX_bit_math_h_l51_c3_edc9_iftrue <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_edc9_iftrue;
     layer0_node3_MUX_bit_math_h_l51_c3_edc9_iffalse <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_edc9_iffalse;
     -- Outputs
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_edc9_return_output := layer0_node3_MUX_bit_math_h_l51_c3_edc9_return_output;

     -- layer0_node16_MUX[bit_math_h_l194_c3_7a7d] LATENCY=0
     -- Inputs
     layer0_node16_MUX_bit_math_h_l194_c3_7a7d_cond <= VAR_layer0_node16_MUX_bit_math_h_l194_c3_7a7d_cond;
     layer0_node16_MUX_bit_math_h_l194_c3_7a7d_iftrue <= VAR_layer0_node16_MUX_bit_math_h_l194_c3_7a7d_iftrue;
     layer0_node16_MUX_bit_math_h_l194_c3_7a7d_iffalse <= VAR_layer0_node16_MUX_bit_math_h_l194_c3_7a7d_iffalse;
     -- Outputs
     VAR_layer0_node16_MUX_bit_math_h_l194_c3_7a7d_return_output := layer0_node16_MUX_bit_math_h_l194_c3_7a7d_return_output;

     -- layer0_node15_MUX[bit_math_h_l183_c3_5274] LATENCY=0
     -- Inputs
     layer0_node15_MUX_bit_math_h_l183_c3_5274_cond <= VAR_layer0_node15_MUX_bit_math_h_l183_c3_5274_cond;
     layer0_node15_MUX_bit_math_h_l183_c3_5274_iftrue <= VAR_layer0_node15_MUX_bit_math_h_l183_c3_5274_iftrue;
     layer0_node15_MUX_bit_math_h_l183_c3_5274_iffalse <= VAR_layer0_node15_MUX_bit_math_h_l183_c3_5274_iffalse;
     -- Outputs
     VAR_layer0_node15_MUX_bit_math_h_l183_c3_5274_return_output := layer0_node15_MUX_bit_math_h_l183_c3_5274_return_output;

     -- layer0_node44_MUX[bit_math_h_l502_c3_15dc] LATENCY=0
     -- Inputs
     layer0_node44_MUX_bit_math_h_l502_c3_15dc_cond <= VAR_layer0_node44_MUX_bit_math_h_l502_c3_15dc_cond;
     layer0_node44_MUX_bit_math_h_l502_c3_15dc_iftrue <= VAR_layer0_node44_MUX_bit_math_h_l502_c3_15dc_iftrue;
     layer0_node44_MUX_bit_math_h_l502_c3_15dc_iffalse <= VAR_layer0_node44_MUX_bit_math_h_l502_c3_15dc_iffalse;
     -- Outputs
     VAR_layer0_node44_MUX_bit_math_h_l502_c3_15dc_return_output := layer0_node44_MUX_bit_math_h_l502_c3_15dc_return_output;

     -- layer0_node20_MUX[bit_math_h_l238_c3_091e] LATENCY=0
     -- Inputs
     layer0_node20_MUX_bit_math_h_l238_c3_091e_cond <= VAR_layer0_node20_MUX_bit_math_h_l238_c3_091e_cond;
     layer0_node20_MUX_bit_math_h_l238_c3_091e_iftrue <= VAR_layer0_node20_MUX_bit_math_h_l238_c3_091e_iftrue;
     layer0_node20_MUX_bit_math_h_l238_c3_091e_iffalse <= VAR_layer0_node20_MUX_bit_math_h_l238_c3_091e_iffalse;
     -- Outputs
     VAR_layer0_node20_MUX_bit_math_h_l238_c3_091e_return_output := layer0_node20_MUX_bit_math_h_l238_c3_091e_return_output;

     -- layer0_node1_MUX[bit_math_h_l29_c3_0e94] LATENCY=0
     -- Inputs
     layer0_node1_MUX_bit_math_h_l29_c3_0e94_cond <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_0e94_cond;
     layer0_node1_MUX_bit_math_h_l29_c3_0e94_iftrue <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_0e94_iftrue;
     layer0_node1_MUX_bit_math_h_l29_c3_0e94_iffalse <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_0e94_iffalse;
     -- Outputs
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_0e94_return_output := layer0_node1_MUX_bit_math_h_l29_c3_0e94_return_output;

     -- layer0_node0_MUX[bit_math_h_l18_c3_ce9b] LATENCY=0
     -- Inputs
     layer0_node0_MUX_bit_math_h_l18_c3_ce9b_cond <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_ce9b_cond;
     layer0_node0_MUX_bit_math_h_l18_c3_ce9b_iftrue <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_ce9b_iftrue;
     layer0_node0_MUX_bit_math_h_l18_c3_ce9b_iffalse <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_ce9b_iffalse;
     -- Outputs
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_ce9b_return_output := layer0_node0_MUX_bit_math_h_l18_c3_ce9b_return_output;

     -- layer0_node37_MUX[bit_math_h_l425_c3_3900] LATENCY=0
     -- Inputs
     layer0_node37_MUX_bit_math_h_l425_c3_3900_cond <= VAR_layer0_node37_MUX_bit_math_h_l425_c3_3900_cond;
     layer0_node37_MUX_bit_math_h_l425_c3_3900_iftrue <= VAR_layer0_node37_MUX_bit_math_h_l425_c3_3900_iftrue;
     layer0_node37_MUX_bit_math_h_l425_c3_3900_iffalse <= VAR_layer0_node37_MUX_bit_math_h_l425_c3_3900_iffalse;
     -- Outputs
     VAR_layer0_node37_MUX_bit_math_h_l425_c3_3900_return_output := layer0_node37_MUX_bit_math_h_l425_c3_3900_return_output;

     -- layer0_node18_MUX[bit_math_h_l216_c3_b8f1] LATENCY=0
     -- Inputs
     layer0_node18_MUX_bit_math_h_l216_c3_b8f1_cond <= VAR_layer0_node18_MUX_bit_math_h_l216_c3_b8f1_cond;
     layer0_node18_MUX_bit_math_h_l216_c3_b8f1_iftrue <= VAR_layer0_node18_MUX_bit_math_h_l216_c3_b8f1_iftrue;
     layer0_node18_MUX_bit_math_h_l216_c3_b8f1_iffalse <= VAR_layer0_node18_MUX_bit_math_h_l216_c3_b8f1_iffalse;
     -- Outputs
     VAR_layer0_node18_MUX_bit_math_h_l216_c3_b8f1_return_output := layer0_node18_MUX_bit_math_h_l216_c3_b8f1_return_output;

     -- layer0_node23_MUX[bit_math_h_l271_c3_0038] LATENCY=0
     -- Inputs
     layer0_node23_MUX_bit_math_h_l271_c3_0038_cond <= VAR_layer0_node23_MUX_bit_math_h_l271_c3_0038_cond;
     layer0_node23_MUX_bit_math_h_l271_c3_0038_iftrue <= VAR_layer0_node23_MUX_bit_math_h_l271_c3_0038_iftrue;
     layer0_node23_MUX_bit_math_h_l271_c3_0038_iffalse <= VAR_layer0_node23_MUX_bit_math_h_l271_c3_0038_iffalse;
     -- Outputs
     VAR_layer0_node23_MUX_bit_math_h_l271_c3_0038_return_output := layer0_node23_MUX_bit_math_h_l271_c3_0038_return_output;

     -- layer0_node56_MUX[bit_math_h_l634_c3_8e72] LATENCY=0
     -- Inputs
     layer0_node56_MUX_bit_math_h_l634_c3_8e72_cond <= VAR_layer0_node56_MUX_bit_math_h_l634_c3_8e72_cond;
     layer0_node56_MUX_bit_math_h_l634_c3_8e72_iftrue <= VAR_layer0_node56_MUX_bit_math_h_l634_c3_8e72_iftrue;
     layer0_node56_MUX_bit_math_h_l634_c3_8e72_iffalse <= VAR_layer0_node56_MUX_bit_math_h_l634_c3_8e72_iffalse;
     -- Outputs
     VAR_layer0_node56_MUX_bit_math_h_l634_c3_8e72_return_output := layer0_node56_MUX_bit_math_h_l634_c3_8e72_return_output;

     -- layer0_node24_MUX[bit_math_h_l282_c3_1d56] LATENCY=0
     -- Inputs
     layer0_node24_MUX_bit_math_h_l282_c3_1d56_cond <= VAR_layer0_node24_MUX_bit_math_h_l282_c3_1d56_cond;
     layer0_node24_MUX_bit_math_h_l282_c3_1d56_iftrue <= VAR_layer0_node24_MUX_bit_math_h_l282_c3_1d56_iftrue;
     layer0_node24_MUX_bit_math_h_l282_c3_1d56_iffalse <= VAR_layer0_node24_MUX_bit_math_h_l282_c3_1d56_iffalse;
     -- Outputs
     VAR_layer0_node24_MUX_bit_math_h_l282_c3_1d56_return_output := layer0_node24_MUX_bit_math_h_l282_c3_1d56_return_output;

     -- layer0_node22_MUX[bit_math_h_l260_c3_db28] LATENCY=0
     -- Inputs
     layer0_node22_MUX_bit_math_h_l260_c3_db28_cond <= VAR_layer0_node22_MUX_bit_math_h_l260_c3_db28_cond;
     layer0_node22_MUX_bit_math_h_l260_c3_db28_iftrue <= VAR_layer0_node22_MUX_bit_math_h_l260_c3_db28_iftrue;
     layer0_node22_MUX_bit_math_h_l260_c3_db28_iffalse <= VAR_layer0_node22_MUX_bit_math_h_l260_c3_db28_iffalse;
     -- Outputs
     VAR_layer0_node22_MUX_bit_math_h_l260_c3_db28_return_output := layer0_node22_MUX_bit_math_h_l260_c3_db28_return_output;

     -- layer0_node30_MUX[bit_math_h_l348_c3_46cf] LATENCY=0
     -- Inputs
     layer0_node30_MUX_bit_math_h_l348_c3_46cf_cond <= VAR_layer0_node30_MUX_bit_math_h_l348_c3_46cf_cond;
     layer0_node30_MUX_bit_math_h_l348_c3_46cf_iftrue <= VAR_layer0_node30_MUX_bit_math_h_l348_c3_46cf_iftrue;
     layer0_node30_MUX_bit_math_h_l348_c3_46cf_iffalse <= VAR_layer0_node30_MUX_bit_math_h_l348_c3_46cf_iffalse;
     -- Outputs
     VAR_layer0_node30_MUX_bit_math_h_l348_c3_46cf_return_output := layer0_node30_MUX_bit_math_h_l348_c3_46cf_return_output;

     -- layer0_node39_MUX[bit_math_h_l447_c3_3acc] LATENCY=0
     -- Inputs
     layer0_node39_MUX_bit_math_h_l447_c3_3acc_cond <= VAR_layer0_node39_MUX_bit_math_h_l447_c3_3acc_cond;
     layer0_node39_MUX_bit_math_h_l447_c3_3acc_iftrue <= VAR_layer0_node39_MUX_bit_math_h_l447_c3_3acc_iftrue;
     layer0_node39_MUX_bit_math_h_l447_c3_3acc_iffalse <= VAR_layer0_node39_MUX_bit_math_h_l447_c3_3acc_iffalse;
     -- Outputs
     VAR_layer0_node39_MUX_bit_math_h_l447_c3_3acc_return_output := layer0_node39_MUX_bit_math_h_l447_c3_3acc_return_output;

     -- layer0_node41_MUX[bit_math_h_l469_c3_2ffe] LATENCY=0
     -- Inputs
     layer0_node41_MUX_bit_math_h_l469_c3_2ffe_cond <= VAR_layer0_node41_MUX_bit_math_h_l469_c3_2ffe_cond;
     layer0_node41_MUX_bit_math_h_l469_c3_2ffe_iftrue <= VAR_layer0_node41_MUX_bit_math_h_l469_c3_2ffe_iftrue;
     layer0_node41_MUX_bit_math_h_l469_c3_2ffe_iffalse <= VAR_layer0_node41_MUX_bit_math_h_l469_c3_2ffe_iffalse;
     -- Outputs
     VAR_layer0_node41_MUX_bit_math_h_l469_c3_2ffe_return_output := layer0_node41_MUX_bit_math_h_l469_c3_2ffe_return_output;

     -- layer0_node38_MUX[bit_math_h_l436_c3_bea2] LATENCY=0
     -- Inputs
     layer0_node38_MUX_bit_math_h_l436_c3_bea2_cond <= VAR_layer0_node38_MUX_bit_math_h_l436_c3_bea2_cond;
     layer0_node38_MUX_bit_math_h_l436_c3_bea2_iftrue <= VAR_layer0_node38_MUX_bit_math_h_l436_c3_bea2_iftrue;
     layer0_node38_MUX_bit_math_h_l436_c3_bea2_iffalse <= VAR_layer0_node38_MUX_bit_math_h_l436_c3_bea2_iffalse;
     -- Outputs
     VAR_layer0_node38_MUX_bit_math_h_l436_c3_bea2_return_output := layer0_node38_MUX_bit_math_h_l436_c3_bea2_return_output;

     -- layer0_node40_MUX[bit_math_h_l458_c3_f867] LATENCY=0
     -- Inputs
     layer0_node40_MUX_bit_math_h_l458_c3_f867_cond <= VAR_layer0_node40_MUX_bit_math_h_l458_c3_f867_cond;
     layer0_node40_MUX_bit_math_h_l458_c3_f867_iftrue <= VAR_layer0_node40_MUX_bit_math_h_l458_c3_f867_iftrue;
     layer0_node40_MUX_bit_math_h_l458_c3_f867_iffalse <= VAR_layer0_node40_MUX_bit_math_h_l458_c3_f867_iffalse;
     -- Outputs
     VAR_layer0_node40_MUX_bit_math_h_l458_c3_f867_return_output := layer0_node40_MUX_bit_math_h_l458_c3_f867_return_output;

     -- Submodule level 2
     VAR_layer1_node0_MUX_bit_math_h_l728_c3_4268_iffalse := VAR_layer0_node0_MUX_bit_math_h_l18_c3_ce9b_return_output;
     VAR_layer1_node5_MUX_bit_math_h_l783_c3_6db3_iffalse := VAR_layer0_node10_MUX_bit_math_h_l128_c3_06f3_return_output;
     VAR_layer1_node5_MUX_bit_math_h_l783_c3_6db3_iftrue := VAR_layer0_node11_MUX_bit_math_h_l139_c3_dbfc_return_output;
     VAR_layer1_node6_MUX_bit_math_h_l794_c3_4c59_iffalse := VAR_layer0_node12_MUX_bit_math_h_l150_c3_6613_return_output;
     VAR_layer1_node6_MUX_bit_math_h_l794_c3_4c59_iftrue := VAR_layer0_node13_MUX_bit_math_h_l161_c3_fd42_return_output;
     VAR_layer1_node7_MUX_bit_math_h_l805_c3_502f_iffalse := VAR_layer0_node14_MUX_bit_math_h_l172_c3_154a_return_output;
     VAR_layer1_node7_MUX_bit_math_h_l805_c3_502f_iftrue := VAR_layer0_node15_MUX_bit_math_h_l183_c3_5274_return_output;
     VAR_layer1_node8_MUX_bit_math_h_l816_c3_1eec_iffalse := VAR_layer0_node16_MUX_bit_math_h_l194_c3_7a7d_return_output;
     VAR_layer1_node8_MUX_bit_math_h_l816_c3_1eec_iftrue := VAR_layer0_node17_MUX_bit_math_h_l205_c3_42ac_return_output;
     VAR_layer1_node9_MUX_bit_math_h_l827_c3_d105_iffalse := VAR_layer0_node18_MUX_bit_math_h_l216_c3_b8f1_return_output;
     VAR_layer1_node9_MUX_bit_math_h_l827_c3_d105_iftrue := VAR_layer0_node19_MUX_bit_math_h_l227_c3_0b12_return_output;
     VAR_layer1_node0_MUX_bit_math_h_l728_c3_4268_iftrue := VAR_layer0_node1_MUX_bit_math_h_l29_c3_0e94_return_output;
     VAR_layer1_node10_MUX_bit_math_h_l838_c3_8a99_iffalse := VAR_layer0_node20_MUX_bit_math_h_l238_c3_091e_return_output;
     VAR_layer1_node10_MUX_bit_math_h_l838_c3_8a99_iftrue := VAR_layer0_node21_MUX_bit_math_h_l249_c3_44d2_return_output;
     VAR_layer1_node11_MUX_bit_math_h_l849_c3_e0a5_iffalse := VAR_layer0_node22_MUX_bit_math_h_l260_c3_db28_return_output;
     VAR_layer1_node11_MUX_bit_math_h_l849_c3_e0a5_iftrue := VAR_layer0_node23_MUX_bit_math_h_l271_c3_0038_return_output;
     VAR_layer1_node12_MUX_bit_math_h_l860_c3_53b9_iffalse := VAR_layer0_node24_MUX_bit_math_h_l282_c3_1d56_return_output;
     VAR_layer1_node12_MUX_bit_math_h_l860_c3_53b9_iftrue := VAR_layer0_node25_MUX_bit_math_h_l293_c3_fa3c_return_output;
     VAR_layer1_node13_MUX_bit_math_h_l871_c3_672a_iffalse := VAR_layer0_node26_MUX_bit_math_h_l304_c3_220e_return_output;
     VAR_layer1_node13_MUX_bit_math_h_l871_c3_672a_iftrue := VAR_layer0_node27_MUX_bit_math_h_l315_c3_37d2_return_output;
     VAR_layer1_node14_MUX_bit_math_h_l882_c3_2725_iffalse := VAR_layer0_node28_MUX_bit_math_h_l326_c3_af14_return_output;
     VAR_layer1_node14_MUX_bit_math_h_l882_c3_2725_iftrue := VAR_layer0_node29_MUX_bit_math_h_l337_c3_d491_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l739_c3_ff28_iffalse := VAR_layer0_node2_MUX_bit_math_h_l40_c3_e2d9_return_output;
     VAR_layer1_node15_MUX_bit_math_h_l893_c3_b457_iffalse := VAR_layer0_node30_MUX_bit_math_h_l348_c3_46cf_return_output;
     VAR_layer1_node15_MUX_bit_math_h_l893_c3_b457_iftrue := VAR_layer0_node31_MUX_bit_math_h_l359_c3_1ee6_return_output;
     VAR_layer1_node16_MUX_bit_math_h_l904_c3_8832_iffalse := VAR_layer0_node32_MUX_bit_math_h_l370_c3_ee39_return_output;
     VAR_layer1_node16_MUX_bit_math_h_l904_c3_8832_iftrue := VAR_layer0_node33_MUX_bit_math_h_l381_c3_f57d_return_output;
     VAR_layer1_node17_MUX_bit_math_h_l915_c3_0128_iffalse := VAR_layer0_node34_MUX_bit_math_h_l392_c3_8d4e_return_output;
     VAR_layer1_node17_MUX_bit_math_h_l915_c3_0128_iftrue := VAR_layer0_node35_MUX_bit_math_h_l403_c3_fa1f_return_output;
     VAR_layer1_node18_MUX_bit_math_h_l926_c3_a8cf_iffalse := VAR_layer0_node36_MUX_bit_math_h_l414_c3_39b4_return_output;
     VAR_layer1_node18_MUX_bit_math_h_l926_c3_a8cf_iftrue := VAR_layer0_node37_MUX_bit_math_h_l425_c3_3900_return_output;
     VAR_layer1_node19_MUX_bit_math_h_l937_c3_3d6b_iffalse := VAR_layer0_node38_MUX_bit_math_h_l436_c3_bea2_return_output;
     VAR_layer1_node19_MUX_bit_math_h_l937_c3_3d6b_iftrue := VAR_layer0_node39_MUX_bit_math_h_l447_c3_3acc_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l739_c3_ff28_iftrue := VAR_layer0_node3_MUX_bit_math_h_l51_c3_edc9_return_output;
     VAR_layer1_node20_MUX_bit_math_h_l948_c3_331f_iffalse := VAR_layer0_node40_MUX_bit_math_h_l458_c3_f867_return_output;
     VAR_layer1_node20_MUX_bit_math_h_l948_c3_331f_iftrue := VAR_layer0_node41_MUX_bit_math_h_l469_c3_2ffe_return_output;
     VAR_layer1_node21_MUX_bit_math_h_l959_c3_32d5_iffalse := VAR_layer0_node42_MUX_bit_math_h_l480_c3_1c62_return_output;
     VAR_layer1_node21_MUX_bit_math_h_l959_c3_32d5_iftrue := VAR_layer0_node43_MUX_bit_math_h_l491_c3_7943_return_output;
     VAR_layer1_node22_MUX_bit_math_h_l970_c3_56f9_iffalse := VAR_layer0_node44_MUX_bit_math_h_l502_c3_15dc_return_output;
     VAR_layer1_node22_MUX_bit_math_h_l970_c3_56f9_iftrue := VAR_layer0_node45_MUX_bit_math_h_l513_c3_d638_return_output;
     VAR_layer1_node23_MUX_bit_math_h_l981_c3_251b_iffalse := VAR_layer0_node46_MUX_bit_math_h_l524_c3_fdc0_return_output;
     VAR_layer1_node23_MUX_bit_math_h_l981_c3_251b_iftrue := VAR_layer0_node47_MUX_bit_math_h_l535_c3_1640_return_output;
     VAR_layer1_node24_MUX_bit_math_h_l992_c3_a508_iffalse := VAR_layer0_node48_MUX_bit_math_h_l546_c3_b0f6_return_output;
     VAR_layer1_node24_MUX_bit_math_h_l992_c3_a508_iftrue := VAR_layer0_node49_MUX_bit_math_h_l557_c3_adcc_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l750_c3_543f_iffalse := VAR_layer0_node4_MUX_bit_math_h_l62_c3_f389_return_output;
     VAR_layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_iffalse := VAR_layer0_node50_MUX_bit_math_h_l568_c3_e90e_return_output;
     VAR_layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_iftrue := VAR_layer0_node51_MUX_bit_math_h_l579_c3_221f_return_output;
     VAR_layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_iffalse := VAR_layer0_node52_MUX_bit_math_h_l590_c3_70e0_return_output;
     VAR_layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_iftrue := VAR_layer0_node53_MUX_bit_math_h_l601_c3_e235_return_output;
     VAR_layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_iffalse := VAR_layer0_node54_MUX_bit_math_h_l612_c3_f982_return_output;
     VAR_layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_iftrue := VAR_layer0_node55_MUX_bit_math_h_l623_c3_bc3d_return_output;
     VAR_layer1_node28_MUX_bit_math_h_l1036_c3_064f_iffalse := VAR_layer0_node56_MUX_bit_math_h_l634_c3_8e72_return_output;
     VAR_layer1_node28_MUX_bit_math_h_l1036_c3_064f_iftrue := VAR_layer0_node57_MUX_bit_math_h_l645_c3_0789_return_output;
     VAR_layer1_node29_MUX_bit_math_h_l1047_c3_e950_iffalse := VAR_layer0_node58_MUX_bit_math_h_l656_c3_d346_return_output;
     VAR_layer1_node29_MUX_bit_math_h_l1047_c3_e950_iftrue := VAR_layer0_node59_MUX_bit_math_h_l667_c3_d31e_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l750_c3_543f_iftrue := VAR_layer0_node5_MUX_bit_math_h_l73_c3_d655_return_output;
     VAR_layer1_node30_MUX_bit_math_h_l1058_c3_fdae_iffalse := VAR_layer0_node60_MUX_bit_math_h_l678_c3_e120_return_output;
     VAR_layer1_node30_MUX_bit_math_h_l1058_c3_fdae_iftrue := VAR_layer0_node61_MUX_bit_math_h_l689_c3_a1a2_return_output;
     VAR_layer1_node31_MUX_bit_math_h_l1069_c3_6030_iffalse := VAR_layer0_node62_MUX_bit_math_h_l700_c3_4595_return_output;
     VAR_layer1_node31_MUX_bit_math_h_l1069_c3_6030_iftrue := VAR_layer0_node63_MUX_bit_math_h_l711_c3_c6ab_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l761_c3_5c18_iffalse := VAR_layer0_node6_MUX_bit_math_h_l84_c3_5cd3_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l761_c3_5c18_iftrue := VAR_layer0_node7_MUX_bit_math_h_l95_c3_5030_return_output;
     VAR_layer1_node4_MUX_bit_math_h_l772_c3_a66b_iffalse := VAR_layer0_node8_MUX_bit_math_h_l106_c3_32cb_return_output;
     VAR_layer1_node4_MUX_bit_math_h_l772_c3_a66b_iftrue := VAR_layer0_node9_MUX_bit_math_h_l117_c3_4b42_return_output;
     -- layer1_node28_MUX[bit_math_h_l1036_c3_064f] LATENCY=0
     -- Inputs
     layer1_node28_MUX_bit_math_h_l1036_c3_064f_cond <= VAR_layer1_node28_MUX_bit_math_h_l1036_c3_064f_cond;
     layer1_node28_MUX_bit_math_h_l1036_c3_064f_iftrue <= VAR_layer1_node28_MUX_bit_math_h_l1036_c3_064f_iftrue;
     layer1_node28_MUX_bit_math_h_l1036_c3_064f_iffalse <= VAR_layer1_node28_MUX_bit_math_h_l1036_c3_064f_iffalse;
     -- Outputs
     VAR_layer1_node28_MUX_bit_math_h_l1036_c3_064f_return_output := layer1_node28_MUX_bit_math_h_l1036_c3_064f_return_output;

     -- layer1_node5_MUX[bit_math_h_l783_c3_6db3] LATENCY=0
     -- Inputs
     layer1_node5_MUX_bit_math_h_l783_c3_6db3_cond <= VAR_layer1_node5_MUX_bit_math_h_l783_c3_6db3_cond;
     layer1_node5_MUX_bit_math_h_l783_c3_6db3_iftrue <= VAR_layer1_node5_MUX_bit_math_h_l783_c3_6db3_iftrue;
     layer1_node5_MUX_bit_math_h_l783_c3_6db3_iffalse <= VAR_layer1_node5_MUX_bit_math_h_l783_c3_6db3_iffalse;
     -- Outputs
     VAR_layer1_node5_MUX_bit_math_h_l783_c3_6db3_return_output := layer1_node5_MUX_bit_math_h_l783_c3_6db3_return_output;

     -- layer1_node30_MUX[bit_math_h_l1058_c3_fdae] LATENCY=0
     -- Inputs
     layer1_node30_MUX_bit_math_h_l1058_c3_fdae_cond <= VAR_layer1_node30_MUX_bit_math_h_l1058_c3_fdae_cond;
     layer1_node30_MUX_bit_math_h_l1058_c3_fdae_iftrue <= VAR_layer1_node30_MUX_bit_math_h_l1058_c3_fdae_iftrue;
     layer1_node30_MUX_bit_math_h_l1058_c3_fdae_iffalse <= VAR_layer1_node30_MUX_bit_math_h_l1058_c3_fdae_iffalse;
     -- Outputs
     VAR_layer1_node30_MUX_bit_math_h_l1058_c3_fdae_return_output := layer1_node30_MUX_bit_math_h_l1058_c3_fdae_return_output;

     -- layer1_node20_MUX[bit_math_h_l948_c3_331f] LATENCY=0
     -- Inputs
     layer1_node20_MUX_bit_math_h_l948_c3_331f_cond <= VAR_layer1_node20_MUX_bit_math_h_l948_c3_331f_cond;
     layer1_node20_MUX_bit_math_h_l948_c3_331f_iftrue <= VAR_layer1_node20_MUX_bit_math_h_l948_c3_331f_iftrue;
     layer1_node20_MUX_bit_math_h_l948_c3_331f_iffalse <= VAR_layer1_node20_MUX_bit_math_h_l948_c3_331f_iffalse;
     -- Outputs
     VAR_layer1_node20_MUX_bit_math_h_l948_c3_331f_return_output := layer1_node20_MUX_bit_math_h_l948_c3_331f_return_output;

     -- layer1_node3_MUX[bit_math_h_l761_c3_5c18] LATENCY=0
     -- Inputs
     layer1_node3_MUX_bit_math_h_l761_c3_5c18_cond <= VAR_layer1_node3_MUX_bit_math_h_l761_c3_5c18_cond;
     layer1_node3_MUX_bit_math_h_l761_c3_5c18_iftrue <= VAR_layer1_node3_MUX_bit_math_h_l761_c3_5c18_iftrue;
     layer1_node3_MUX_bit_math_h_l761_c3_5c18_iffalse <= VAR_layer1_node3_MUX_bit_math_h_l761_c3_5c18_iffalse;
     -- Outputs
     VAR_layer1_node3_MUX_bit_math_h_l761_c3_5c18_return_output := layer1_node3_MUX_bit_math_h_l761_c3_5c18_return_output;

     -- layer1_node31_MUX[bit_math_h_l1069_c3_6030] LATENCY=0
     -- Inputs
     layer1_node31_MUX_bit_math_h_l1069_c3_6030_cond <= VAR_layer1_node31_MUX_bit_math_h_l1069_c3_6030_cond;
     layer1_node31_MUX_bit_math_h_l1069_c3_6030_iftrue <= VAR_layer1_node31_MUX_bit_math_h_l1069_c3_6030_iftrue;
     layer1_node31_MUX_bit_math_h_l1069_c3_6030_iffalse <= VAR_layer1_node31_MUX_bit_math_h_l1069_c3_6030_iffalse;
     -- Outputs
     VAR_layer1_node31_MUX_bit_math_h_l1069_c3_6030_return_output := layer1_node31_MUX_bit_math_h_l1069_c3_6030_return_output;

     -- layer1_node24_MUX[bit_math_h_l992_c3_a508] LATENCY=0
     -- Inputs
     layer1_node24_MUX_bit_math_h_l992_c3_a508_cond <= VAR_layer1_node24_MUX_bit_math_h_l992_c3_a508_cond;
     layer1_node24_MUX_bit_math_h_l992_c3_a508_iftrue <= VAR_layer1_node24_MUX_bit_math_h_l992_c3_a508_iftrue;
     layer1_node24_MUX_bit_math_h_l992_c3_a508_iffalse <= VAR_layer1_node24_MUX_bit_math_h_l992_c3_a508_iffalse;
     -- Outputs
     VAR_layer1_node24_MUX_bit_math_h_l992_c3_a508_return_output := layer1_node24_MUX_bit_math_h_l992_c3_a508_return_output;

     -- layer1_node8_MUX[bit_math_h_l816_c3_1eec] LATENCY=0
     -- Inputs
     layer1_node8_MUX_bit_math_h_l816_c3_1eec_cond <= VAR_layer1_node8_MUX_bit_math_h_l816_c3_1eec_cond;
     layer1_node8_MUX_bit_math_h_l816_c3_1eec_iftrue <= VAR_layer1_node8_MUX_bit_math_h_l816_c3_1eec_iftrue;
     layer1_node8_MUX_bit_math_h_l816_c3_1eec_iffalse <= VAR_layer1_node8_MUX_bit_math_h_l816_c3_1eec_iffalse;
     -- Outputs
     VAR_layer1_node8_MUX_bit_math_h_l816_c3_1eec_return_output := layer1_node8_MUX_bit_math_h_l816_c3_1eec_return_output;

     -- layer1_node29_MUX[bit_math_h_l1047_c3_e950] LATENCY=0
     -- Inputs
     layer1_node29_MUX_bit_math_h_l1047_c3_e950_cond <= VAR_layer1_node29_MUX_bit_math_h_l1047_c3_e950_cond;
     layer1_node29_MUX_bit_math_h_l1047_c3_e950_iftrue <= VAR_layer1_node29_MUX_bit_math_h_l1047_c3_e950_iftrue;
     layer1_node29_MUX_bit_math_h_l1047_c3_e950_iffalse <= VAR_layer1_node29_MUX_bit_math_h_l1047_c3_e950_iffalse;
     -- Outputs
     VAR_layer1_node29_MUX_bit_math_h_l1047_c3_e950_return_output := layer1_node29_MUX_bit_math_h_l1047_c3_e950_return_output;

     -- layer1_node14_MUX[bit_math_h_l882_c3_2725] LATENCY=0
     -- Inputs
     layer1_node14_MUX_bit_math_h_l882_c3_2725_cond <= VAR_layer1_node14_MUX_bit_math_h_l882_c3_2725_cond;
     layer1_node14_MUX_bit_math_h_l882_c3_2725_iftrue <= VAR_layer1_node14_MUX_bit_math_h_l882_c3_2725_iftrue;
     layer1_node14_MUX_bit_math_h_l882_c3_2725_iffalse <= VAR_layer1_node14_MUX_bit_math_h_l882_c3_2725_iffalse;
     -- Outputs
     VAR_layer1_node14_MUX_bit_math_h_l882_c3_2725_return_output := layer1_node14_MUX_bit_math_h_l882_c3_2725_return_output;

     -- layer1_node4_MUX[bit_math_h_l772_c3_a66b] LATENCY=0
     -- Inputs
     layer1_node4_MUX_bit_math_h_l772_c3_a66b_cond <= VAR_layer1_node4_MUX_bit_math_h_l772_c3_a66b_cond;
     layer1_node4_MUX_bit_math_h_l772_c3_a66b_iftrue <= VAR_layer1_node4_MUX_bit_math_h_l772_c3_a66b_iftrue;
     layer1_node4_MUX_bit_math_h_l772_c3_a66b_iffalse <= VAR_layer1_node4_MUX_bit_math_h_l772_c3_a66b_iffalse;
     -- Outputs
     VAR_layer1_node4_MUX_bit_math_h_l772_c3_a66b_return_output := layer1_node4_MUX_bit_math_h_l772_c3_a66b_return_output;

     -- layer1_node25_MUX[bit_math_h_l1003_c3_6bb3] LATENCY=0
     -- Inputs
     layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_cond <= VAR_layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_cond;
     layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_iftrue <= VAR_layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_iftrue;
     layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_iffalse <= VAR_layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_iffalse;
     -- Outputs
     VAR_layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_return_output := layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_return_output;

     -- layer1_node26_MUX[bit_math_h_l1014_c3_5bdb] LATENCY=0
     -- Inputs
     layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_cond <= VAR_layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_cond;
     layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_iftrue <= VAR_layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_iftrue;
     layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_iffalse <= VAR_layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_iffalse;
     -- Outputs
     VAR_layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_return_output := layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_return_output;

     -- layer1_node18_MUX[bit_math_h_l926_c3_a8cf] LATENCY=0
     -- Inputs
     layer1_node18_MUX_bit_math_h_l926_c3_a8cf_cond <= VAR_layer1_node18_MUX_bit_math_h_l926_c3_a8cf_cond;
     layer1_node18_MUX_bit_math_h_l926_c3_a8cf_iftrue <= VAR_layer1_node18_MUX_bit_math_h_l926_c3_a8cf_iftrue;
     layer1_node18_MUX_bit_math_h_l926_c3_a8cf_iffalse <= VAR_layer1_node18_MUX_bit_math_h_l926_c3_a8cf_iffalse;
     -- Outputs
     VAR_layer1_node18_MUX_bit_math_h_l926_c3_a8cf_return_output := layer1_node18_MUX_bit_math_h_l926_c3_a8cf_return_output;

     -- layer1_node21_MUX[bit_math_h_l959_c3_32d5] LATENCY=0
     -- Inputs
     layer1_node21_MUX_bit_math_h_l959_c3_32d5_cond <= VAR_layer1_node21_MUX_bit_math_h_l959_c3_32d5_cond;
     layer1_node21_MUX_bit_math_h_l959_c3_32d5_iftrue <= VAR_layer1_node21_MUX_bit_math_h_l959_c3_32d5_iftrue;
     layer1_node21_MUX_bit_math_h_l959_c3_32d5_iffalse <= VAR_layer1_node21_MUX_bit_math_h_l959_c3_32d5_iffalse;
     -- Outputs
     VAR_layer1_node21_MUX_bit_math_h_l959_c3_32d5_return_output := layer1_node21_MUX_bit_math_h_l959_c3_32d5_return_output;

     -- layer1_node11_MUX[bit_math_h_l849_c3_e0a5] LATENCY=0
     -- Inputs
     layer1_node11_MUX_bit_math_h_l849_c3_e0a5_cond <= VAR_layer1_node11_MUX_bit_math_h_l849_c3_e0a5_cond;
     layer1_node11_MUX_bit_math_h_l849_c3_e0a5_iftrue <= VAR_layer1_node11_MUX_bit_math_h_l849_c3_e0a5_iftrue;
     layer1_node11_MUX_bit_math_h_l849_c3_e0a5_iffalse <= VAR_layer1_node11_MUX_bit_math_h_l849_c3_e0a5_iffalse;
     -- Outputs
     VAR_layer1_node11_MUX_bit_math_h_l849_c3_e0a5_return_output := layer1_node11_MUX_bit_math_h_l849_c3_e0a5_return_output;

     -- layer1_node22_MUX[bit_math_h_l970_c3_56f9] LATENCY=0
     -- Inputs
     layer1_node22_MUX_bit_math_h_l970_c3_56f9_cond <= VAR_layer1_node22_MUX_bit_math_h_l970_c3_56f9_cond;
     layer1_node22_MUX_bit_math_h_l970_c3_56f9_iftrue <= VAR_layer1_node22_MUX_bit_math_h_l970_c3_56f9_iftrue;
     layer1_node22_MUX_bit_math_h_l970_c3_56f9_iffalse <= VAR_layer1_node22_MUX_bit_math_h_l970_c3_56f9_iffalse;
     -- Outputs
     VAR_layer1_node22_MUX_bit_math_h_l970_c3_56f9_return_output := layer1_node22_MUX_bit_math_h_l970_c3_56f9_return_output;

     -- layer1_node7_MUX[bit_math_h_l805_c3_502f] LATENCY=0
     -- Inputs
     layer1_node7_MUX_bit_math_h_l805_c3_502f_cond <= VAR_layer1_node7_MUX_bit_math_h_l805_c3_502f_cond;
     layer1_node7_MUX_bit_math_h_l805_c3_502f_iftrue <= VAR_layer1_node7_MUX_bit_math_h_l805_c3_502f_iftrue;
     layer1_node7_MUX_bit_math_h_l805_c3_502f_iffalse <= VAR_layer1_node7_MUX_bit_math_h_l805_c3_502f_iffalse;
     -- Outputs
     VAR_layer1_node7_MUX_bit_math_h_l805_c3_502f_return_output := layer1_node7_MUX_bit_math_h_l805_c3_502f_return_output;

     -- layer1_node0_MUX[bit_math_h_l728_c3_4268] LATENCY=0
     -- Inputs
     layer1_node0_MUX_bit_math_h_l728_c3_4268_cond <= VAR_layer1_node0_MUX_bit_math_h_l728_c3_4268_cond;
     layer1_node0_MUX_bit_math_h_l728_c3_4268_iftrue <= VAR_layer1_node0_MUX_bit_math_h_l728_c3_4268_iftrue;
     layer1_node0_MUX_bit_math_h_l728_c3_4268_iffalse <= VAR_layer1_node0_MUX_bit_math_h_l728_c3_4268_iffalse;
     -- Outputs
     VAR_layer1_node0_MUX_bit_math_h_l728_c3_4268_return_output := layer1_node0_MUX_bit_math_h_l728_c3_4268_return_output;

     -- layer1_node12_MUX[bit_math_h_l860_c3_53b9] LATENCY=0
     -- Inputs
     layer1_node12_MUX_bit_math_h_l860_c3_53b9_cond <= VAR_layer1_node12_MUX_bit_math_h_l860_c3_53b9_cond;
     layer1_node12_MUX_bit_math_h_l860_c3_53b9_iftrue <= VAR_layer1_node12_MUX_bit_math_h_l860_c3_53b9_iftrue;
     layer1_node12_MUX_bit_math_h_l860_c3_53b9_iffalse <= VAR_layer1_node12_MUX_bit_math_h_l860_c3_53b9_iffalse;
     -- Outputs
     VAR_layer1_node12_MUX_bit_math_h_l860_c3_53b9_return_output := layer1_node12_MUX_bit_math_h_l860_c3_53b9_return_output;

     -- layer1_node15_MUX[bit_math_h_l893_c3_b457] LATENCY=0
     -- Inputs
     layer1_node15_MUX_bit_math_h_l893_c3_b457_cond <= VAR_layer1_node15_MUX_bit_math_h_l893_c3_b457_cond;
     layer1_node15_MUX_bit_math_h_l893_c3_b457_iftrue <= VAR_layer1_node15_MUX_bit_math_h_l893_c3_b457_iftrue;
     layer1_node15_MUX_bit_math_h_l893_c3_b457_iffalse <= VAR_layer1_node15_MUX_bit_math_h_l893_c3_b457_iffalse;
     -- Outputs
     VAR_layer1_node15_MUX_bit_math_h_l893_c3_b457_return_output := layer1_node15_MUX_bit_math_h_l893_c3_b457_return_output;

     -- layer1_node16_MUX[bit_math_h_l904_c3_8832] LATENCY=0
     -- Inputs
     layer1_node16_MUX_bit_math_h_l904_c3_8832_cond <= VAR_layer1_node16_MUX_bit_math_h_l904_c3_8832_cond;
     layer1_node16_MUX_bit_math_h_l904_c3_8832_iftrue <= VAR_layer1_node16_MUX_bit_math_h_l904_c3_8832_iftrue;
     layer1_node16_MUX_bit_math_h_l904_c3_8832_iffalse <= VAR_layer1_node16_MUX_bit_math_h_l904_c3_8832_iffalse;
     -- Outputs
     VAR_layer1_node16_MUX_bit_math_h_l904_c3_8832_return_output := layer1_node16_MUX_bit_math_h_l904_c3_8832_return_output;

     -- layer1_node27_MUX[bit_math_h_l1025_c3_a0dc] LATENCY=0
     -- Inputs
     layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_cond <= VAR_layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_cond;
     layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_iftrue <= VAR_layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_iftrue;
     layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_iffalse <= VAR_layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_iffalse;
     -- Outputs
     VAR_layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_return_output := layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_return_output;

     -- layer1_node9_MUX[bit_math_h_l827_c3_d105] LATENCY=0
     -- Inputs
     layer1_node9_MUX_bit_math_h_l827_c3_d105_cond <= VAR_layer1_node9_MUX_bit_math_h_l827_c3_d105_cond;
     layer1_node9_MUX_bit_math_h_l827_c3_d105_iftrue <= VAR_layer1_node9_MUX_bit_math_h_l827_c3_d105_iftrue;
     layer1_node9_MUX_bit_math_h_l827_c3_d105_iffalse <= VAR_layer1_node9_MUX_bit_math_h_l827_c3_d105_iffalse;
     -- Outputs
     VAR_layer1_node9_MUX_bit_math_h_l827_c3_d105_return_output := layer1_node9_MUX_bit_math_h_l827_c3_d105_return_output;

     -- layer1_node13_MUX[bit_math_h_l871_c3_672a] LATENCY=0
     -- Inputs
     layer1_node13_MUX_bit_math_h_l871_c3_672a_cond <= VAR_layer1_node13_MUX_bit_math_h_l871_c3_672a_cond;
     layer1_node13_MUX_bit_math_h_l871_c3_672a_iftrue <= VAR_layer1_node13_MUX_bit_math_h_l871_c3_672a_iftrue;
     layer1_node13_MUX_bit_math_h_l871_c3_672a_iffalse <= VAR_layer1_node13_MUX_bit_math_h_l871_c3_672a_iffalse;
     -- Outputs
     VAR_layer1_node13_MUX_bit_math_h_l871_c3_672a_return_output := layer1_node13_MUX_bit_math_h_l871_c3_672a_return_output;

     -- layer1_node10_MUX[bit_math_h_l838_c3_8a99] LATENCY=0
     -- Inputs
     layer1_node10_MUX_bit_math_h_l838_c3_8a99_cond <= VAR_layer1_node10_MUX_bit_math_h_l838_c3_8a99_cond;
     layer1_node10_MUX_bit_math_h_l838_c3_8a99_iftrue <= VAR_layer1_node10_MUX_bit_math_h_l838_c3_8a99_iftrue;
     layer1_node10_MUX_bit_math_h_l838_c3_8a99_iffalse <= VAR_layer1_node10_MUX_bit_math_h_l838_c3_8a99_iffalse;
     -- Outputs
     VAR_layer1_node10_MUX_bit_math_h_l838_c3_8a99_return_output := layer1_node10_MUX_bit_math_h_l838_c3_8a99_return_output;

     -- layer1_node2_MUX[bit_math_h_l750_c3_543f] LATENCY=0
     -- Inputs
     layer1_node2_MUX_bit_math_h_l750_c3_543f_cond <= VAR_layer1_node2_MUX_bit_math_h_l750_c3_543f_cond;
     layer1_node2_MUX_bit_math_h_l750_c3_543f_iftrue <= VAR_layer1_node2_MUX_bit_math_h_l750_c3_543f_iftrue;
     layer1_node2_MUX_bit_math_h_l750_c3_543f_iffalse <= VAR_layer1_node2_MUX_bit_math_h_l750_c3_543f_iffalse;
     -- Outputs
     VAR_layer1_node2_MUX_bit_math_h_l750_c3_543f_return_output := layer1_node2_MUX_bit_math_h_l750_c3_543f_return_output;

     -- layer1_node19_MUX[bit_math_h_l937_c3_3d6b] LATENCY=0
     -- Inputs
     layer1_node19_MUX_bit_math_h_l937_c3_3d6b_cond <= VAR_layer1_node19_MUX_bit_math_h_l937_c3_3d6b_cond;
     layer1_node19_MUX_bit_math_h_l937_c3_3d6b_iftrue <= VAR_layer1_node19_MUX_bit_math_h_l937_c3_3d6b_iftrue;
     layer1_node19_MUX_bit_math_h_l937_c3_3d6b_iffalse <= VAR_layer1_node19_MUX_bit_math_h_l937_c3_3d6b_iffalse;
     -- Outputs
     VAR_layer1_node19_MUX_bit_math_h_l937_c3_3d6b_return_output := layer1_node19_MUX_bit_math_h_l937_c3_3d6b_return_output;

     -- layer1_node1_MUX[bit_math_h_l739_c3_ff28] LATENCY=0
     -- Inputs
     layer1_node1_MUX_bit_math_h_l739_c3_ff28_cond <= VAR_layer1_node1_MUX_bit_math_h_l739_c3_ff28_cond;
     layer1_node1_MUX_bit_math_h_l739_c3_ff28_iftrue <= VAR_layer1_node1_MUX_bit_math_h_l739_c3_ff28_iftrue;
     layer1_node1_MUX_bit_math_h_l739_c3_ff28_iffalse <= VAR_layer1_node1_MUX_bit_math_h_l739_c3_ff28_iffalse;
     -- Outputs
     VAR_layer1_node1_MUX_bit_math_h_l739_c3_ff28_return_output := layer1_node1_MUX_bit_math_h_l739_c3_ff28_return_output;

     -- layer1_node17_MUX[bit_math_h_l915_c3_0128] LATENCY=0
     -- Inputs
     layer1_node17_MUX_bit_math_h_l915_c3_0128_cond <= VAR_layer1_node17_MUX_bit_math_h_l915_c3_0128_cond;
     layer1_node17_MUX_bit_math_h_l915_c3_0128_iftrue <= VAR_layer1_node17_MUX_bit_math_h_l915_c3_0128_iftrue;
     layer1_node17_MUX_bit_math_h_l915_c3_0128_iffalse <= VAR_layer1_node17_MUX_bit_math_h_l915_c3_0128_iffalse;
     -- Outputs
     VAR_layer1_node17_MUX_bit_math_h_l915_c3_0128_return_output := layer1_node17_MUX_bit_math_h_l915_c3_0128_return_output;

     -- layer1_node6_MUX[bit_math_h_l794_c3_4c59] LATENCY=0
     -- Inputs
     layer1_node6_MUX_bit_math_h_l794_c3_4c59_cond <= VAR_layer1_node6_MUX_bit_math_h_l794_c3_4c59_cond;
     layer1_node6_MUX_bit_math_h_l794_c3_4c59_iftrue <= VAR_layer1_node6_MUX_bit_math_h_l794_c3_4c59_iftrue;
     layer1_node6_MUX_bit_math_h_l794_c3_4c59_iffalse <= VAR_layer1_node6_MUX_bit_math_h_l794_c3_4c59_iffalse;
     -- Outputs
     VAR_layer1_node6_MUX_bit_math_h_l794_c3_4c59_return_output := layer1_node6_MUX_bit_math_h_l794_c3_4c59_return_output;

     -- layer1_node23_MUX[bit_math_h_l981_c3_251b] LATENCY=0
     -- Inputs
     layer1_node23_MUX_bit_math_h_l981_c3_251b_cond <= VAR_layer1_node23_MUX_bit_math_h_l981_c3_251b_cond;
     layer1_node23_MUX_bit_math_h_l981_c3_251b_iftrue <= VAR_layer1_node23_MUX_bit_math_h_l981_c3_251b_iftrue;
     layer1_node23_MUX_bit_math_h_l981_c3_251b_iffalse <= VAR_layer1_node23_MUX_bit_math_h_l981_c3_251b_iffalse;
     -- Outputs
     VAR_layer1_node23_MUX_bit_math_h_l981_c3_251b_return_output := layer1_node23_MUX_bit_math_h_l981_c3_251b_return_output;

     -- Submodule level 3
     VAR_layer2_node0_MUX_bit_math_h_l1086_c3_122d_iffalse := VAR_layer1_node0_MUX_bit_math_h_l728_c3_4268_return_output;
     VAR_layer2_node5_MUX_bit_math_h_l1141_c3_1425_iffalse := VAR_layer1_node10_MUX_bit_math_h_l838_c3_8a99_return_output;
     VAR_layer2_node5_MUX_bit_math_h_l1141_c3_1425_iftrue := VAR_layer1_node11_MUX_bit_math_h_l849_c3_e0a5_return_output;
     VAR_layer2_node6_MUX_bit_math_h_l1152_c3_008a_iffalse := VAR_layer1_node12_MUX_bit_math_h_l860_c3_53b9_return_output;
     VAR_layer2_node6_MUX_bit_math_h_l1152_c3_008a_iftrue := VAR_layer1_node13_MUX_bit_math_h_l871_c3_672a_return_output;
     VAR_layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_iffalse := VAR_layer1_node14_MUX_bit_math_h_l882_c3_2725_return_output;
     VAR_layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_iftrue := VAR_layer1_node15_MUX_bit_math_h_l893_c3_b457_return_output;
     VAR_layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_iffalse := VAR_layer1_node16_MUX_bit_math_h_l904_c3_8832_return_output;
     VAR_layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_iftrue := VAR_layer1_node17_MUX_bit_math_h_l915_c3_0128_return_output;
     VAR_layer2_node9_MUX_bit_math_h_l1185_c3_98c3_iffalse := VAR_layer1_node18_MUX_bit_math_h_l926_c3_a8cf_return_output;
     VAR_layer2_node9_MUX_bit_math_h_l1185_c3_98c3_iftrue := VAR_layer1_node19_MUX_bit_math_h_l937_c3_3d6b_return_output;
     VAR_layer2_node0_MUX_bit_math_h_l1086_c3_122d_iftrue := VAR_layer1_node1_MUX_bit_math_h_l739_c3_ff28_return_output;
     VAR_layer2_node10_MUX_bit_math_h_l1196_c3_1666_iffalse := VAR_layer1_node20_MUX_bit_math_h_l948_c3_331f_return_output;
     VAR_layer2_node10_MUX_bit_math_h_l1196_c3_1666_iftrue := VAR_layer1_node21_MUX_bit_math_h_l959_c3_32d5_return_output;
     VAR_layer2_node11_MUX_bit_math_h_l1207_c3_b8de_iffalse := VAR_layer1_node22_MUX_bit_math_h_l970_c3_56f9_return_output;
     VAR_layer2_node11_MUX_bit_math_h_l1207_c3_b8de_iftrue := VAR_layer1_node23_MUX_bit_math_h_l981_c3_251b_return_output;
     VAR_layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_iffalse := VAR_layer1_node24_MUX_bit_math_h_l992_c3_a508_return_output;
     VAR_layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_iftrue := VAR_layer1_node25_MUX_bit_math_h_l1003_c3_6bb3_return_output;
     VAR_layer2_node13_MUX_bit_math_h_l1229_c3_d585_iffalse := VAR_layer1_node26_MUX_bit_math_h_l1014_c3_5bdb_return_output;
     VAR_layer2_node13_MUX_bit_math_h_l1229_c3_d585_iftrue := VAR_layer1_node27_MUX_bit_math_h_l1025_c3_a0dc_return_output;
     VAR_layer2_node14_MUX_bit_math_h_l1240_c3_beb5_iffalse := VAR_layer1_node28_MUX_bit_math_h_l1036_c3_064f_return_output;
     VAR_layer2_node14_MUX_bit_math_h_l1240_c3_beb5_iftrue := VAR_layer1_node29_MUX_bit_math_h_l1047_c3_e950_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_iffalse := VAR_layer1_node2_MUX_bit_math_h_l750_c3_543f_return_output;
     VAR_layer2_node15_MUX_bit_math_h_l1251_c3_7550_iffalse := VAR_layer1_node30_MUX_bit_math_h_l1058_c3_fdae_return_output;
     VAR_layer2_node15_MUX_bit_math_h_l1251_c3_7550_iftrue := VAR_layer1_node31_MUX_bit_math_h_l1069_c3_6030_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_iftrue := VAR_layer1_node3_MUX_bit_math_h_l761_c3_5c18_return_output;
     VAR_layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_iffalse := VAR_layer1_node4_MUX_bit_math_h_l772_c3_a66b_return_output;
     VAR_layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_iftrue := VAR_layer1_node5_MUX_bit_math_h_l783_c3_6db3_return_output;
     VAR_layer2_node3_MUX_bit_math_h_l1119_c3_946d_iffalse := VAR_layer1_node6_MUX_bit_math_h_l794_c3_4c59_return_output;
     VAR_layer2_node3_MUX_bit_math_h_l1119_c3_946d_iftrue := VAR_layer1_node7_MUX_bit_math_h_l805_c3_502f_return_output;
     VAR_layer2_node4_MUX_bit_math_h_l1130_c3_1f93_iffalse := VAR_layer1_node8_MUX_bit_math_h_l816_c3_1eec_return_output;
     VAR_layer2_node4_MUX_bit_math_h_l1130_c3_1f93_iftrue := VAR_layer1_node9_MUX_bit_math_h_l827_c3_d105_return_output;
     -- layer2_node11_MUX[bit_math_h_l1207_c3_b8de] LATENCY=0
     -- Inputs
     layer2_node11_MUX_bit_math_h_l1207_c3_b8de_cond <= VAR_layer2_node11_MUX_bit_math_h_l1207_c3_b8de_cond;
     layer2_node11_MUX_bit_math_h_l1207_c3_b8de_iftrue <= VAR_layer2_node11_MUX_bit_math_h_l1207_c3_b8de_iftrue;
     layer2_node11_MUX_bit_math_h_l1207_c3_b8de_iffalse <= VAR_layer2_node11_MUX_bit_math_h_l1207_c3_b8de_iffalse;
     -- Outputs
     VAR_layer2_node11_MUX_bit_math_h_l1207_c3_b8de_return_output := layer2_node11_MUX_bit_math_h_l1207_c3_b8de_return_output;

     -- layer2_node2_MUX[bit_math_h_l1108_c3_b1b3] LATENCY=0
     -- Inputs
     layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_cond <= VAR_layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_cond;
     layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_iftrue <= VAR_layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_iftrue;
     layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_iffalse <= VAR_layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_iffalse;
     -- Outputs
     VAR_layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_return_output := layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_return_output;

     -- layer2_node1_MUX[bit_math_h_l1097_c3_fcc7] LATENCY=0
     -- Inputs
     layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_cond <= VAR_layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_cond;
     layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_iftrue <= VAR_layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_iftrue;
     layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_iffalse <= VAR_layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_iffalse;
     -- Outputs
     VAR_layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_return_output := layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_return_output;

     -- layer2_node14_MUX[bit_math_h_l1240_c3_beb5] LATENCY=0
     -- Inputs
     layer2_node14_MUX_bit_math_h_l1240_c3_beb5_cond <= VAR_layer2_node14_MUX_bit_math_h_l1240_c3_beb5_cond;
     layer2_node14_MUX_bit_math_h_l1240_c3_beb5_iftrue <= VAR_layer2_node14_MUX_bit_math_h_l1240_c3_beb5_iftrue;
     layer2_node14_MUX_bit_math_h_l1240_c3_beb5_iffalse <= VAR_layer2_node14_MUX_bit_math_h_l1240_c3_beb5_iffalse;
     -- Outputs
     VAR_layer2_node14_MUX_bit_math_h_l1240_c3_beb5_return_output := layer2_node14_MUX_bit_math_h_l1240_c3_beb5_return_output;

     -- layer2_node15_MUX[bit_math_h_l1251_c3_7550] LATENCY=0
     -- Inputs
     layer2_node15_MUX_bit_math_h_l1251_c3_7550_cond <= VAR_layer2_node15_MUX_bit_math_h_l1251_c3_7550_cond;
     layer2_node15_MUX_bit_math_h_l1251_c3_7550_iftrue <= VAR_layer2_node15_MUX_bit_math_h_l1251_c3_7550_iftrue;
     layer2_node15_MUX_bit_math_h_l1251_c3_7550_iffalse <= VAR_layer2_node15_MUX_bit_math_h_l1251_c3_7550_iffalse;
     -- Outputs
     VAR_layer2_node15_MUX_bit_math_h_l1251_c3_7550_return_output := layer2_node15_MUX_bit_math_h_l1251_c3_7550_return_output;

     -- layer2_node0_MUX[bit_math_h_l1086_c3_122d] LATENCY=0
     -- Inputs
     layer2_node0_MUX_bit_math_h_l1086_c3_122d_cond <= VAR_layer2_node0_MUX_bit_math_h_l1086_c3_122d_cond;
     layer2_node0_MUX_bit_math_h_l1086_c3_122d_iftrue <= VAR_layer2_node0_MUX_bit_math_h_l1086_c3_122d_iftrue;
     layer2_node0_MUX_bit_math_h_l1086_c3_122d_iffalse <= VAR_layer2_node0_MUX_bit_math_h_l1086_c3_122d_iffalse;
     -- Outputs
     VAR_layer2_node0_MUX_bit_math_h_l1086_c3_122d_return_output := layer2_node0_MUX_bit_math_h_l1086_c3_122d_return_output;

     -- layer2_node10_MUX[bit_math_h_l1196_c3_1666] LATENCY=0
     -- Inputs
     layer2_node10_MUX_bit_math_h_l1196_c3_1666_cond <= VAR_layer2_node10_MUX_bit_math_h_l1196_c3_1666_cond;
     layer2_node10_MUX_bit_math_h_l1196_c3_1666_iftrue <= VAR_layer2_node10_MUX_bit_math_h_l1196_c3_1666_iftrue;
     layer2_node10_MUX_bit_math_h_l1196_c3_1666_iffalse <= VAR_layer2_node10_MUX_bit_math_h_l1196_c3_1666_iffalse;
     -- Outputs
     VAR_layer2_node10_MUX_bit_math_h_l1196_c3_1666_return_output := layer2_node10_MUX_bit_math_h_l1196_c3_1666_return_output;

     -- layer2_node7_MUX[bit_math_h_l1163_c3_5ba0] LATENCY=0
     -- Inputs
     layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_cond <= VAR_layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_cond;
     layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_iftrue <= VAR_layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_iftrue;
     layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_iffalse <= VAR_layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_iffalse;
     -- Outputs
     VAR_layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_return_output := layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_return_output;

     -- layer2_node13_MUX[bit_math_h_l1229_c3_d585] LATENCY=0
     -- Inputs
     layer2_node13_MUX_bit_math_h_l1229_c3_d585_cond <= VAR_layer2_node13_MUX_bit_math_h_l1229_c3_d585_cond;
     layer2_node13_MUX_bit_math_h_l1229_c3_d585_iftrue <= VAR_layer2_node13_MUX_bit_math_h_l1229_c3_d585_iftrue;
     layer2_node13_MUX_bit_math_h_l1229_c3_d585_iffalse <= VAR_layer2_node13_MUX_bit_math_h_l1229_c3_d585_iffalse;
     -- Outputs
     VAR_layer2_node13_MUX_bit_math_h_l1229_c3_d585_return_output := layer2_node13_MUX_bit_math_h_l1229_c3_d585_return_output;

     -- layer2_node4_MUX[bit_math_h_l1130_c3_1f93] LATENCY=0
     -- Inputs
     layer2_node4_MUX_bit_math_h_l1130_c3_1f93_cond <= VAR_layer2_node4_MUX_bit_math_h_l1130_c3_1f93_cond;
     layer2_node4_MUX_bit_math_h_l1130_c3_1f93_iftrue <= VAR_layer2_node4_MUX_bit_math_h_l1130_c3_1f93_iftrue;
     layer2_node4_MUX_bit_math_h_l1130_c3_1f93_iffalse <= VAR_layer2_node4_MUX_bit_math_h_l1130_c3_1f93_iffalse;
     -- Outputs
     VAR_layer2_node4_MUX_bit_math_h_l1130_c3_1f93_return_output := layer2_node4_MUX_bit_math_h_l1130_c3_1f93_return_output;

     -- layer2_node5_MUX[bit_math_h_l1141_c3_1425] LATENCY=0
     -- Inputs
     layer2_node5_MUX_bit_math_h_l1141_c3_1425_cond <= VAR_layer2_node5_MUX_bit_math_h_l1141_c3_1425_cond;
     layer2_node5_MUX_bit_math_h_l1141_c3_1425_iftrue <= VAR_layer2_node5_MUX_bit_math_h_l1141_c3_1425_iftrue;
     layer2_node5_MUX_bit_math_h_l1141_c3_1425_iffalse <= VAR_layer2_node5_MUX_bit_math_h_l1141_c3_1425_iffalse;
     -- Outputs
     VAR_layer2_node5_MUX_bit_math_h_l1141_c3_1425_return_output := layer2_node5_MUX_bit_math_h_l1141_c3_1425_return_output;

     -- layer2_node6_MUX[bit_math_h_l1152_c3_008a] LATENCY=0
     -- Inputs
     layer2_node6_MUX_bit_math_h_l1152_c3_008a_cond <= VAR_layer2_node6_MUX_bit_math_h_l1152_c3_008a_cond;
     layer2_node6_MUX_bit_math_h_l1152_c3_008a_iftrue <= VAR_layer2_node6_MUX_bit_math_h_l1152_c3_008a_iftrue;
     layer2_node6_MUX_bit_math_h_l1152_c3_008a_iffalse <= VAR_layer2_node6_MUX_bit_math_h_l1152_c3_008a_iffalse;
     -- Outputs
     VAR_layer2_node6_MUX_bit_math_h_l1152_c3_008a_return_output := layer2_node6_MUX_bit_math_h_l1152_c3_008a_return_output;

     -- layer2_node8_MUX[bit_math_h_l1174_c3_f1cf] LATENCY=0
     -- Inputs
     layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_cond <= VAR_layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_cond;
     layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_iftrue <= VAR_layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_iftrue;
     layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_iffalse <= VAR_layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_iffalse;
     -- Outputs
     VAR_layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_return_output := layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_return_output;

     -- layer2_node9_MUX[bit_math_h_l1185_c3_98c3] LATENCY=0
     -- Inputs
     layer2_node9_MUX_bit_math_h_l1185_c3_98c3_cond <= VAR_layer2_node9_MUX_bit_math_h_l1185_c3_98c3_cond;
     layer2_node9_MUX_bit_math_h_l1185_c3_98c3_iftrue <= VAR_layer2_node9_MUX_bit_math_h_l1185_c3_98c3_iftrue;
     layer2_node9_MUX_bit_math_h_l1185_c3_98c3_iffalse <= VAR_layer2_node9_MUX_bit_math_h_l1185_c3_98c3_iffalse;
     -- Outputs
     VAR_layer2_node9_MUX_bit_math_h_l1185_c3_98c3_return_output := layer2_node9_MUX_bit_math_h_l1185_c3_98c3_return_output;

     -- layer2_node3_MUX[bit_math_h_l1119_c3_946d] LATENCY=0
     -- Inputs
     layer2_node3_MUX_bit_math_h_l1119_c3_946d_cond <= VAR_layer2_node3_MUX_bit_math_h_l1119_c3_946d_cond;
     layer2_node3_MUX_bit_math_h_l1119_c3_946d_iftrue <= VAR_layer2_node3_MUX_bit_math_h_l1119_c3_946d_iftrue;
     layer2_node3_MUX_bit_math_h_l1119_c3_946d_iffalse <= VAR_layer2_node3_MUX_bit_math_h_l1119_c3_946d_iffalse;
     -- Outputs
     VAR_layer2_node3_MUX_bit_math_h_l1119_c3_946d_return_output := layer2_node3_MUX_bit_math_h_l1119_c3_946d_return_output;

     -- layer2_node12_MUX[bit_math_h_l1218_c3_d8dc] LATENCY=0
     -- Inputs
     layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_cond <= VAR_layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_cond;
     layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_iftrue <= VAR_layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_iftrue;
     layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_iffalse <= VAR_layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_iffalse;
     -- Outputs
     VAR_layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_return_output := layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_return_output;

     -- Submodule level 4
     VAR_layer3_node0_MUX_bit_math_h_l1268_c3_302d_iffalse := VAR_layer2_node0_MUX_bit_math_h_l1086_c3_122d_return_output;
     VAR_layer3_node5_MUX_bit_math_h_l1323_c3_57ee_iffalse := VAR_layer2_node10_MUX_bit_math_h_l1196_c3_1666_return_output;
     VAR_layer3_node5_MUX_bit_math_h_l1323_c3_57ee_iftrue := VAR_layer2_node11_MUX_bit_math_h_l1207_c3_b8de_return_output;
     VAR_layer3_node6_MUX_bit_math_h_l1334_c3_f24c_iffalse := VAR_layer2_node12_MUX_bit_math_h_l1218_c3_d8dc_return_output;
     VAR_layer3_node6_MUX_bit_math_h_l1334_c3_f24c_iftrue := VAR_layer2_node13_MUX_bit_math_h_l1229_c3_d585_return_output;
     VAR_layer3_node7_MUX_bit_math_h_l1345_c3_c68c_iffalse := VAR_layer2_node14_MUX_bit_math_h_l1240_c3_beb5_return_output;
     VAR_layer3_node7_MUX_bit_math_h_l1345_c3_c68c_iftrue := VAR_layer2_node15_MUX_bit_math_h_l1251_c3_7550_return_output;
     VAR_layer3_node0_MUX_bit_math_h_l1268_c3_302d_iftrue := VAR_layer2_node1_MUX_bit_math_h_l1097_c3_fcc7_return_output;
     VAR_layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_iffalse := VAR_layer2_node2_MUX_bit_math_h_l1108_c3_b1b3_return_output;
     VAR_layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_iftrue := VAR_layer2_node3_MUX_bit_math_h_l1119_c3_946d_return_output;
     VAR_layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_iffalse := VAR_layer2_node4_MUX_bit_math_h_l1130_c3_1f93_return_output;
     VAR_layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_iftrue := VAR_layer2_node5_MUX_bit_math_h_l1141_c3_1425_return_output;
     VAR_layer3_node3_MUX_bit_math_h_l1301_c3_84c3_iffalse := VAR_layer2_node6_MUX_bit_math_h_l1152_c3_008a_return_output;
     VAR_layer3_node3_MUX_bit_math_h_l1301_c3_84c3_iftrue := VAR_layer2_node7_MUX_bit_math_h_l1163_c3_5ba0_return_output;
     VAR_layer3_node4_MUX_bit_math_h_l1312_c3_8c96_iffalse := VAR_layer2_node8_MUX_bit_math_h_l1174_c3_f1cf_return_output;
     VAR_layer3_node4_MUX_bit_math_h_l1312_c3_8c96_iftrue := VAR_layer2_node9_MUX_bit_math_h_l1185_c3_98c3_return_output;
     -- layer3_node0_MUX[bit_math_h_l1268_c3_302d] LATENCY=0
     -- Inputs
     layer3_node0_MUX_bit_math_h_l1268_c3_302d_cond <= VAR_layer3_node0_MUX_bit_math_h_l1268_c3_302d_cond;
     layer3_node0_MUX_bit_math_h_l1268_c3_302d_iftrue <= VAR_layer3_node0_MUX_bit_math_h_l1268_c3_302d_iftrue;
     layer3_node0_MUX_bit_math_h_l1268_c3_302d_iffalse <= VAR_layer3_node0_MUX_bit_math_h_l1268_c3_302d_iffalse;
     -- Outputs
     VAR_layer3_node0_MUX_bit_math_h_l1268_c3_302d_return_output := layer3_node0_MUX_bit_math_h_l1268_c3_302d_return_output;

     -- layer3_node6_MUX[bit_math_h_l1334_c3_f24c] LATENCY=0
     -- Inputs
     layer3_node6_MUX_bit_math_h_l1334_c3_f24c_cond <= VAR_layer3_node6_MUX_bit_math_h_l1334_c3_f24c_cond;
     layer3_node6_MUX_bit_math_h_l1334_c3_f24c_iftrue <= VAR_layer3_node6_MUX_bit_math_h_l1334_c3_f24c_iftrue;
     layer3_node6_MUX_bit_math_h_l1334_c3_f24c_iffalse <= VAR_layer3_node6_MUX_bit_math_h_l1334_c3_f24c_iffalse;
     -- Outputs
     VAR_layer3_node6_MUX_bit_math_h_l1334_c3_f24c_return_output := layer3_node6_MUX_bit_math_h_l1334_c3_f24c_return_output;

     -- layer3_node5_MUX[bit_math_h_l1323_c3_57ee] LATENCY=0
     -- Inputs
     layer3_node5_MUX_bit_math_h_l1323_c3_57ee_cond <= VAR_layer3_node5_MUX_bit_math_h_l1323_c3_57ee_cond;
     layer3_node5_MUX_bit_math_h_l1323_c3_57ee_iftrue <= VAR_layer3_node5_MUX_bit_math_h_l1323_c3_57ee_iftrue;
     layer3_node5_MUX_bit_math_h_l1323_c3_57ee_iffalse <= VAR_layer3_node5_MUX_bit_math_h_l1323_c3_57ee_iffalse;
     -- Outputs
     VAR_layer3_node5_MUX_bit_math_h_l1323_c3_57ee_return_output := layer3_node5_MUX_bit_math_h_l1323_c3_57ee_return_output;

     -- layer3_node7_MUX[bit_math_h_l1345_c3_c68c] LATENCY=0
     -- Inputs
     layer3_node7_MUX_bit_math_h_l1345_c3_c68c_cond <= VAR_layer3_node7_MUX_bit_math_h_l1345_c3_c68c_cond;
     layer3_node7_MUX_bit_math_h_l1345_c3_c68c_iftrue <= VAR_layer3_node7_MUX_bit_math_h_l1345_c3_c68c_iftrue;
     layer3_node7_MUX_bit_math_h_l1345_c3_c68c_iffalse <= VAR_layer3_node7_MUX_bit_math_h_l1345_c3_c68c_iffalse;
     -- Outputs
     VAR_layer3_node7_MUX_bit_math_h_l1345_c3_c68c_return_output := layer3_node7_MUX_bit_math_h_l1345_c3_c68c_return_output;

     -- layer3_node3_MUX[bit_math_h_l1301_c3_84c3] LATENCY=0
     -- Inputs
     layer3_node3_MUX_bit_math_h_l1301_c3_84c3_cond <= VAR_layer3_node3_MUX_bit_math_h_l1301_c3_84c3_cond;
     layer3_node3_MUX_bit_math_h_l1301_c3_84c3_iftrue <= VAR_layer3_node3_MUX_bit_math_h_l1301_c3_84c3_iftrue;
     layer3_node3_MUX_bit_math_h_l1301_c3_84c3_iffalse <= VAR_layer3_node3_MUX_bit_math_h_l1301_c3_84c3_iffalse;
     -- Outputs
     VAR_layer3_node3_MUX_bit_math_h_l1301_c3_84c3_return_output := layer3_node3_MUX_bit_math_h_l1301_c3_84c3_return_output;

     -- layer3_node1_MUX[bit_math_h_l1279_c3_fd3b] LATENCY=0
     -- Inputs
     layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_cond <= VAR_layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_cond;
     layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_iftrue <= VAR_layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_iftrue;
     layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_iffalse <= VAR_layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_iffalse;
     -- Outputs
     VAR_layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_return_output := layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_return_output;

     -- layer3_node4_MUX[bit_math_h_l1312_c3_8c96] LATENCY=0
     -- Inputs
     layer3_node4_MUX_bit_math_h_l1312_c3_8c96_cond <= VAR_layer3_node4_MUX_bit_math_h_l1312_c3_8c96_cond;
     layer3_node4_MUX_bit_math_h_l1312_c3_8c96_iftrue <= VAR_layer3_node4_MUX_bit_math_h_l1312_c3_8c96_iftrue;
     layer3_node4_MUX_bit_math_h_l1312_c3_8c96_iffalse <= VAR_layer3_node4_MUX_bit_math_h_l1312_c3_8c96_iffalse;
     -- Outputs
     VAR_layer3_node4_MUX_bit_math_h_l1312_c3_8c96_return_output := layer3_node4_MUX_bit_math_h_l1312_c3_8c96_return_output;

     -- layer3_node2_MUX[bit_math_h_l1290_c3_5e3f] LATENCY=0
     -- Inputs
     layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_cond <= VAR_layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_cond;
     layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_iftrue <= VAR_layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_iftrue;
     layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_iffalse <= VAR_layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_iffalse;
     -- Outputs
     VAR_layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_return_output := layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_return_output;

     -- Submodule level 5
     VAR_layer4_node0_MUX_bit_math_h_l1362_c3_a122_iffalse := VAR_layer3_node0_MUX_bit_math_h_l1268_c3_302d_return_output;
     VAR_layer4_node0_MUX_bit_math_h_l1362_c3_a122_iftrue := VAR_layer3_node1_MUX_bit_math_h_l1279_c3_fd3b_return_output;
     VAR_layer4_node1_MUX_bit_math_h_l1373_c3_c86f_iffalse := VAR_layer3_node2_MUX_bit_math_h_l1290_c3_5e3f_return_output;
     VAR_layer4_node1_MUX_bit_math_h_l1373_c3_c86f_iftrue := VAR_layer3_node3_MUX_bit_math_h_l1301_c3_84c3_return_output;
     VAR_layer4_node2_MUX_bit_math_h_l1384_c3_76f0_iffalse := VAR_layer3_node4_MUX_bit_math_h_l1312_c3_8c96_return_output;
     VAR_layer4_node2_MUX_bit_math_h_l1384_c3_76f0_iftrue := VAR_layer3_node5_MUX_bit_math_h_l1323_c3_57ee_return_output;
     VAR_layer4_node3_MUX_bit_math_h_l1395_c3_5649_iffalse := VAR_layer3_node6_MUX_bit_math_h_l1334_c3_f24c_return_output;
     VAR_layer4_node3_MUX_bit_math_h_l1395_c3_5649_iftrue := VAR_layer3_node7_MUX_bit_math_h_l1345_c3_c68c_return_output;
     -- layer4_node0_MUX[bit_math_h_l1362_c3_a122] LATENCY=0
     -- Inputs
     layer4_node0_MUX_bit_math_h_l1362_c3_a122_cond <= VAR_layer4_node0_MUX_bit_math_h_l1362_c3_a122_cond;
     layer4_node0_MUX_bit_math_h_l1362_c3_a122_iftrue <= VAR_layer4_node0_MUX_bit_math_h_l1362_c3_a122_iftrue;
     layer4_node0_MUX_bit_math_h_l1362_c3_a122_iffalse <= VAR_layer4_node0_MUX_bit_math_h_l1362_c3_a122_iffalse;
     -- Outputs
     VAR_layer4_node0_MUX_bit_math_h_l1362_c3_a122_return_output := layer4_node0_MUX_bit_math_h_l1362_c3_a122_return_output;

     -- layer4_node3_MUX[bit_math_h_l1395_c3_5649] LATENCY=0
     -- Inputs
     layer4_node3_MUX_bit_math_h_l1395_c3_5649_cond <= VAR_layer4_node3_MUX_bit_math_h_l1395_c3_5649_cond;
     layer4_node3_MUX_bit_math_h_l1395_c3_5649_iftrue <= VAR_layer4_node3_MUX_bit_math_h_l1395_c3_5649_iftrue;
     layer4_node3_MUX_bit_math_h_l1395_c3_5649_iffalse <= VAR_layer4_node3_MUX_bit_math_h_l1395_c3_5649_iffalse;
     -- Outputs
     VAR_layer4_node3_MUX_bit_math_h_l1395_c3_5649_return_output := layer4_node3_MUX_bit_math_h_l1395_c3_5649_return_output;

     -- layer4_node1_MUX[bit_math_h_l1373_c3_c86f] LATENCY=0
     -- Inputs
     layer4_node1_MUX_bit_math_h_l1373_c3_c86f_cond <= VAR_layer4_node1_MUX_bit_math_h_l1373_c3_c86f_cond;
     layer4_node1_MUX_bit_math_h_l1373_c3_c86f_iftrue <= VAR_layer4_node1_MUX_bit_math_h_l1373_c3_c86f_iftrue;
     layer4_node1_MUX_bit_math_h_l1373_c3_c86f_iffalse <= VAR_layer4_node1_MUX_bit_math_h_l1373_c3_c86f_iffalse;
     -- Outputs
     VAR_layer4_node1_MUX_bit_math_h_l1373_c3_c86f_return_output := layer4_node1_MUX_bit_math_h_l1373_c3_c86f_return_output;

     -- layer4_node2_MUX[bit_math_h_l1384_c3_76f0] LATENCY=0
     -- Inputs
     layer4_node2_MUX_bit_math_h_l1384_c3_76f0_cond <= VAR_layer4_node2_MUX_bit_math_h_l1384_c3_76f0_cond;
     layer4_node2_MUX_bit_math_h_l1384_c3_76f0_iftrue <= VAR_layer4_node2_MUX_bit_math_h_l1384_c3_76f0_iftrue;
     layer4_node2_MUX_bit_math_h_l1384_c3_76f0_iffalse <= VAR_layer4_node2_MUX_bit_math_h_l1384_c3_76f0_iffalse;
     -- Outputs
     VAR_layer4_node2_MUX_bit_math_h_l1384_c3_76f0_return_output := layer4_node2_MUX_bit_math_h_l1384_c3_76f0_return_output;

     -- Submodule level 6
     VAR_layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_iffalse := VAR_layer4_node0_MUX_bit_math_h_l1362_c3_a122_return_output;
     VAR_layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_iftrue := VAR_layer4_node1_MUX_bit_math_h_l1373_c3_c86f_return_output;
     VAR_layer5_node1_MUX_bit_math_h_l1423_c3_d92a_iffalse := VAR_layer4_node2_MUX_bit_math_h_l1384_c3_76f0_return_output;
     VAR_layer5_node1_MUX_bit_math_h_l1423_c3_d92a_iftrue := VAR_layer4_node3_MUX_bit_math_h_l1395_c3_5649_return_output;
     -- layer5_node0_MUX[bit_math_h_l1412_c3_c6a2] LATENCY=0
     -- Inputs
     layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_cond <= VAR_layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_cond;
     layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_iftrue <= VAR_layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_iftrue;
     layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_iffalse <= VAR_layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_iffalse;
     -- Outputs
     VAR_layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_return_output := layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_return_output;

     -- layer5_node1_MUX[bit_math_h_l1423_c3_d92a] LATENCY=0
     -- Inputs
     layer5_node1_MUX_bit_math_h_l1423_c3_d92a_cond <= VAR_layer5_node1_MUX_bit_math_h_l1423_c3_d92a_cond;
     layer5_node1_MUX_bit_math_h_l1423_c3_d92a_iftrue <= VAR_layer5_node1_MUX_bit_math_h_l1423_c3_d92a_iftrue;
     layer5_node1_MUX_bit_math_h_l1423_c3_d92a_iffalse <= VAR_layer5_node1_MUX_bit_math_h_l1423_c3_d92a_iffalse;
     -- Outputs
     VAR_layer5_node1_MUX_bit_math_h_l1423_c3_d92a_return_output := layer5_node1_MUX_bit_math_h_l1423_c3_d92a_return_output;

     -- Submodule level 7
     VAR_layer6_node0_MUX_bit_math_h_l1440_c3_43c9_iffalse := VAR_layer5_node0_MUX_bit_math_h_l1412_c3_c6a2_return_output;
     VAR_layer6_node0_MUX_bit_math_h_l1440_c3_43c9_iftrue := VAR_layer5_node1_MUX_bit_math_h_l1423_c3_d92a_return_output;
     -- layer6_node0_MUX[bit_math_h_l1440_c3_43c9] LATENCY=0
     -- Inputs
     layer6_node0_MUX_bit_math_h_l1440_c3_43c9_cond <= VAR_layer6_node0_MUX_bit_math_h_l1440_c3_43c9_cond;
     layer6_node0_MUX_bit_math_h_l1440_c3_43c9_iftrue <= VAR_layer6_node0_MUX_bit_math_h_l1440_c3_43c9_iftrue;
     layer6_node0_MUX_bit_math_h_l1440_c3_43c9_iffalse <= VAR_layer6_node0_MUX_bit_math_h_l1440_c3_43c9_iffalse;
     -- Outputs
     VAR_layer6_node0_MUX_bit_math_h_l1440_c3_43c9_return_output := layer6_node0_MUX_bit_math_h_l1440_c3_43c9_return_output;

     -- Submodule level 8
     VAR_return_output := VAR_layer6_node0_MUX_bit_math_h_l1440_c3_43c9_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
