-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity sft_0CLK_46cced44 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sft_0CLK_46cced44;
architecture arch of sft_0CLK_46cced44 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2213_c6_5770]
signal BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2213_c2_3307]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2213_c2_3307]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2213_c2_3307]
signal result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2213_c2_3307]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2213_c2_3307]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2213_c2_3307]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2213_c2_3307]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2213_c2_3307]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2213_c2_3307]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2213_c2_3307]
signal tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2213_c2_3307]
signal n8_MUX_uxn_opcodes_h_l2213_c2_3307_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2213_c2_3307]
signal t8_MUX_uxn_opcodes_h_l2213_c2_3307_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2226_c11_4e1f]
signal BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2226_c7_41d8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2226_c7_41d8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2226_c7_41d8]
signal result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2226_c7_41d8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2226_c7_41d8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2226_c7_41d8]
signal tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2226_c7_41d8]
signal n8_MUX_uxn_opcodes_h_l2226_c7_41d8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2226_c7_41d8]
signal t8_MUX_uxn_opcodes_h_l2226_c7_41d8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2229_c11_05f4]
signal BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2229_c7_ad46]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2229_c7_ad46]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2229_c7_ad46]
signal result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2229_c7_ad46]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2229_c7_ad46]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2229_c7_ad46]
signal tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2229_c7_ad46]
signal n8_MUX_uxn_opcodes_h_l2229_c7_ad46_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2229_c7_ad46]
signal t8_MUX_uxn_opcodes_h_l2229_c7_ad46_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2231_c30_952c]
signal sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2233_c11_bfc9]
signal BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2233_c7_a443]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2233_c7_a443]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2233_c7_a443]
signal result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2233_c7_a443]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2233_c7_a443]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2233_c7_a443]
signal tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2233_c7_a443]
signal n8_MUX_uxn_opcodes_h_l2233_c7_a443_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2233_c7_a443_return_output : unsigned(7 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l2236_c18_aea4]
signal BIN_OP_AND_uxn_opcodes_h_l2236_c18_aea4_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2236_c18_aea4_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2236_c18_aea4_return_output : unsigned(7 downto 0);

-- BIN_OP_SR[uxn_opcodes_h_l2236_c11_d643]
signal BIN_OP_SR_uxn_opcodes_h_l2236_c11_d643_left : unsigned(7 downto 0);
signal BIN_OP_SR_uxn_opcodes_h_l2236_c11_d643_right : unsigned(7 downto 0);
signal BIN_OP_SR_uxn_opcodes_h_l2236_c11_d643_return_output : unsigned(7 downto 0);

-- CONST_SR_4[uxn_opcodes_h_l2236_c34_0d96]
signal CONST_SR_4_uxn_opcodes_h_l2236_c34_0d96_x : unsigned(7 downto 0);
signal CONST_SR_4_uxn_opcodes_h_l2236_c34_0d96_return_output : unsigned(7 downto 0);

-- BIN_OP_SL[uxn_opcodes_h_l2236_c11_ba52]
signal BIN_OP_SL_uxn_opcodes_h_l2236_c11_ba52_left : unsigned(7 downto 0);
signal BIN_OP_SL_uxn_opcodes_h_l2236_c11_ba52_right : unsigned(7 downto 0);
signal BIN_OP_SL_uxn_opcodes_h_l2236_c11_ba52_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_pc_updated := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.is_ram_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;
      base.is_stack_index_flipped := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770
BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_left,
BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_right,
BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307
result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307
result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307
result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_cond,
result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307
result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2213_c2_3307
tmp8_MUX_uxn_opcodes_h_l2213_c2_3307 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_cond,
tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue,
tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse,
tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_return_output);

-- n8_MUX_uxn_opcodes_h_l2213_c2_3307
n8_MUX_uxn_opcodes_h_l2213_c2_3307 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2213_c2_3307_cond,
n8_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue,
n8_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse,
n8_MUX_uxn_opcodes_h_l2213_c2_3307_return_output);

-- t8_MUX_uxn_opcodes_h_l2213_c2_3307
t8_MUX_uxn_opcodes_h_l2213_c2_3307 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2213_c2_3307_cond,
t8_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue,
t8_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse,
t8_MUX_uxn_opcodes_h_l2213_c2_3307_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f
BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_left,
BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_right,
BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8
result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8
result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8
result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_cond,
result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8
result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8
tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_cond,
tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue,
tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse,
tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output);

-- n8_MUX_uxn_opcodes_h_l2226_c7_41d8
n8_MUX_uxn_opcodes_h_l2226_c7_41d8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2226_c7_41d8_cond,
n8_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue,
n8_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse,
n8_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output);

-- t8_MUX_uxn_opcodes_h_l2226_c7_41d8
t8_MUX_uxn_opcodes_h_l2226_c7_41d8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2226_c7_41d8_cond,
t8_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue,
t8_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse,
t8_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4
BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_left,
BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_right,
BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46
result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46
result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46
result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_cond,
result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46
result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46
tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_cond,
tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue,
tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse,
tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output);

-- n8_MUX_uxn_opcodes_h_l2229_c7_ad46
n8_MUX_uxn_opcodes_h_l2229_c7_ad46 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2229_c7_ad46_cond,
n8_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue,
n8_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse,
n8_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output);

-- t8_MUX_uxn_opcodes_h_l2229_c7_ad46
t8_MUX_uxn_opcodes_h_l2229_c7_ad46 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2229_c7_ad46_cond,
t8_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue,
t8_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse,
t8_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2231_c30_952c
sp_relative_shift_uxn_opcodes_h_l2231_c30_952c : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_ins,
sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_x,
sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_y,
sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9
BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_left,
BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_right,
BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443
result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443
result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443
result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_cond,
result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443
result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2233_c7_a443
tmp8_MUX_uxn_opcodes_h_l2233_c7_a443 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_cond,
tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue,
tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse,
tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_return_output);

-- n8_MUX_uxn_opcodes_h_l2233_c7_a443
n8_MUX_uxn_opcodes_h_l2233_c7_a443 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2233_c7_a443_cond,
n8_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue,
n8_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse,
n8_MUX_uxn_opcodes_h_l2233_c7_a443_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l2236_c18_aea4
BIN_OP_AND_uxn_opcodes_h_l2236_c18_aea4 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l2236_c18_aea4_left,
BIN_OP_AND_uxn_opcodes_h_l2236_c18_aea4_right,
BIN_OP_AND_uxn_opcodes_h_l2236_c18_aea4_return_output);

-- BIN_OP_SR_uxn_opcodes_h_l2236_c11_d643
BIN_OP_SR_uxn_opcodes_h_l2236_c11_d643 : entity work.BIN_OP_SR_uint8_t_uint8_t_0CLK_25d197a7 port map (
BIN_OP_SR_uxn_opcodes_h_l2236_c11_d643_left,
BIN_OP_SR_uxn_opcodes_h_l2236_c11_d643_right,
BIN_OP_SR_uxn_opcodes_h_l2236_c11_d643_return_output);

-- CONST_SR_4_uxn_opcodes_h_l2236_c34_0d96
CONST_SR_4_uxn_opcodes_h_l2236_c34_0d96 : entity work.CONST_SR_4_uint8_t_0CLK_de264c78 port map (
CONST_SR_4_uxn_opcodes_h_l2236_c34_0d96_x,
CONST_SR_4_uxn_opcodes_h_l2236_c34_0d96_return_output);

-- BIN_OP_SL_uxn_opcodes_h_l2236_c11_ba52
BIN_OP_SL_uxn_opcodes_h_l2236_c11_ba52 : entity work.BIN_OP_SL_uint8_t_uint8_t_0CLK_10d8c973 port map (
BIN_OP_SL_uxn_opcodes_h_l2236_c11_ba52_left,
BIN_OP_SL_uxn_opcodes_h_l2236_c11_ba52_right,
BIN_OP_SL_uxn_opcodes_h_l2236_c11_ba52_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_return_output,
 tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_return_output,
 n8_MUX_uxn_opcodes_h_l2213_c2_3307_return_output,
 t8_MUX_uxn_opcodes_h_l2213_c2_3307_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output,
 tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output,
 n8_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output,
 t8_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output,
 tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output,
 n8_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output,
 t8_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output,
 sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_return_output,
 tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_return_output,
 n8_MUX_uxn_opcodes_h_l2233_c7_a443_return_output,
 BIN_OP_AND_uxn_opcodes_h_l2236_c18_aea4_return_output,
 BIN_OP_SR_uxn_opcodes_h_l2236_c11_d643_return_output,
 CONST_SR_4_uxn_opcodes_h_l2236_c34_0d96_return_output,
 BIN_OP_SL_uxn_opcodes_h_l2236_c11_ba52_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2218_c3_2ceb : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2223_c3_6335 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2213_c2_3307_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2213_c2_3307_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2213_c2_3307_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2227_c3_33d0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2226_c7_41d8_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2226_c7_41d8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2233_c7_a443_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2229_c7_ad46_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2229_c7_ad46_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2235_c3_9c6b : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2238_c3_d78a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2233_c7_a443_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_d643_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_aea4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_aea4_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_aea4_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_d643_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_d643_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_ba52_left : unsigned(7 downto 0);
 variable VAR_CONST_SR_4_uxn_opcodes_h_l2236_c34_0d96_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_ba52_right : unsigned(7 downto 0);
 variable VAR_CONST_SR_4_uxn_opcodes_h_l2236_c34_0d96_x : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_ba52_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2229_l2213_l2233_l2226_DUPLICATE_3cd1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2233_l2226_DUPLICATE_26e7_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2229_l2233_l2226_DUPLICATE_9412_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2229_l2233_l2226_DUPLICATE_feb3_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2229_l2233_DUPLICATE_0d56_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l2243_l2209_DUPLICATE_685e_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_aea4_right := to_unsigned(15, 8);
     VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2218_c3_2ceb := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2218_c3_2ceb;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2227_c3_33d0 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2227_c3_33d0;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2235_c3_9c6b := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2235_c3_9c6b;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2238_c3_d78a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2238_c3_d78a;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2223_c3_6335 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2223_c3_6335;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_left := VAR_phase;
     VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_d643_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_aea4_left := t8;
     VAR_CONST_SR_4_uxn_opcodes_h_l2236_c34_0d96_x := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse := tmp8;
     -- sp_relative_shift[uxn_opcodes_h_l2231_c30_952c] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_ins;
     sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_x;
     sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_return_output := sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2229_l2213_l2233_l2226_DUPLICATE_3cd1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2229_l2213_l2233_l2226_DUPLICATE_3cd1_return_output := result.u8_value;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2213_c2_3307] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2213_c2_3307_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2229_l2233_l2226_DUPLICATE_9412 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2229_l2233_l2226_DUPLICATE_9412_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2229_c11_05f4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_left;
     BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_return_output := BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2226_c11_4e1f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_return_output;

     -- CONST_SR_4[uxn_opcodes_h_l2236_c34_0d96] LATENCY=0
     -- Inputs
     CONST_SR_4_uxn_opcodes_h_l2236_c34_0d96_x <= VAR_CONST_SR_4_uxn_opcodes_h_l2236_c34_0d96_x;
     -- Outputs
     VAR_CONST_SR_4_uxn_opcodes_h_l2236_c34_0d96_return_output := CONST_SR_4_uxn_opcodes_h_l2236_c34_0d96_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2213_c2_3307] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2213_c2_3307_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l2233_c11_bfc9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_left;
     BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_return_output := BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2229_l2233_l2226_DUPLICATE_feb3 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2229_l2233_l2226_DUPLICATE_feb3_return_output := result.is_opc_done;

     -- BIN_OP_AND[uxn_opcodes_h_l2236_c18_aea4] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l2236_c18_aea4_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_aea4_left;
     BIN_OP_AND_uxn_opcodes_h_l2236_c18_aea4_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_aea4_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_aea4_return_output := BIN_OP_AND_uxn_opcodes_h_l2236_c18_aea4_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2233_l2226_DUPLICATE_26e7 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2233_l2226_DUPLICATE_26e7_return_output := result.sp_relative_shift;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2213_c2_3307] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2213_c2_3307_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2229_l2233_DUPLICATE_0d56 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2229_l2233_DUPLICATE_0d56_return_output := result.stack_address_sp_offset;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2213_c2_3307] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2213_c2_3307_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2213_c6_5770] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_left;
     BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_return_output := BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_return_output;

     -- Submodule level 1
     VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_d643_right := VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_aea4_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2213_c2_3307_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2213_c2_3307_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_5770_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2226_c7_41d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2226_c7_41d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_4e1f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2229_c7_ad46_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2229_c7_ad46_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_05f4_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2233_c7_a443_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_bfc9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2233_l2226_DUPLICATE_26e7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2233_l2226_DUPLICATE_26e7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2229_l2233_l2226_DUPLICATE_feb3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2229_l2233_l2226_DUPLICATE_feb3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2229_l2233_l2226_DUPLICATE_feb3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2229_l2233_l2226_DUPLICATE_9412_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2229_l2233_l2226_DUPLICATE_9412_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2229_l2233_l2226_DUPLICATE_9412_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2229_l2233_DUPLICATE_0d56_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2229_l2233_DUPLICATE_0d56_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2229_l2213_l2233_l2226_DUPLICATE_3cd1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2229_l2213_l2233_l2226_DUPLICATE_3cd1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2229_l2213_l2233_l2226_DUPLICATE_3cd1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2229_l2213_l2233_l2226_DUPLICATE_3cd1_return_output;
     VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_ba52_right := VAR_CONST_SR_4_uxn_opcodes_h_l2236_c34_0d96_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2213_c2_3307_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2213_c2_3307_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2213_c2_3307_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2213_c2_3307_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_952c_return_output;
     -- result_is_vram_write_MUX[uxn_opcodes_h_l2213_c2_3307] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2213_c2_3307] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2233_c7_a443] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2213_c2_3307] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2233_c7_a443] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2233_c7_a443] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2213_c2_3307] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_return_output;

     -- BIN_OP_SR[uxn_opcodes_h_l2236_c11_d643] LATENCY=0
     -- Inputs
     BIN_OP_SR_uxn_opcodes_h_l2236_c11_d643_left <= VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_d643_left;
     BIN_OP_SR_uxn_opcodes_h_l2236_c11_d643_right <= VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_d643_right;
     -- Outputs
     VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_d643_return_output := BIN_OP_SR_uxn_opcodes_h_l2236_c11_d643_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2233_c7_a443] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_return_output;

     -- n8_MUX[uxn_opcodes_h_l2233_c7_a443] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2233_c7_a443_cond <= VAR_n8_MUX_uxn_opcodes_h_l2233_c7_a443_cond;
     n8_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue;
     n8_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2233_c7_a443_return_output := n8_MUX_uxn_opcodes_h_l2233_c7_a443_return_output;

     -- t8_MUX[uxn_opcodes_h_l2229_c7_ad46] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2229_c7_ad46_cond <= VAR_t8_MUX_uxn_opcodes_h_l2229_c7_ad46_cond;
     t8_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue;
     t8_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output := t8_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output;

     -- Submodule level 2
     VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_ba52_left := VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_d643_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2233_c7_a443_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_a443_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_a443_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_a443_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_a443_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2229_c7_ad46] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2229_c7_ad46] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output;

     -- t8_MUX[uxn_opcodes_h_l2226_c7_41d8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2226_c7_41d8_cond <= VAR_t8_MUX_uxn_opcodes_h_l2226_c7_41d8_cond;
     t8_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue;
     t8_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output := t8_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output;

     -- BIN_OP_SL[uxn_opcodes_h_l2236_c11_ba52] LATENCY=0
     -- Inputs
     BIN_OP_SL_uxn_opcodes_h_l2236_c11_ba52_left <= VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_ba52_left;
     BIN_OP_SL_uxn_opcodes_h_l2236_c11_ba52_right <= VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_ba52_right;
     -- Outputs
     VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_ba52_return_output := BIN_OP_SL_uxn_opcodes_h_l2236_c11_ba52_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2229_c7_ad46] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output;

     -- n8_MUX[uxn_opcodes_h_l2229_c7_ad46] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2229_c7_ad46_cond <= VAR_n8_MUX_uxn_opcodes_h_l2229_c7_ad46_cond;
     n8_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue;
     n8_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output := n8_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2229_c7_ad46] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output;

     -- Submodule level 3
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue := VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_ba52_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue := VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_ba52_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output;
     -- t8_MUX[uxn_opcodes_h_l2213_c2_3307] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2213_c2_3307_cond <= VAR_t8_MUX_uxn_opcodes_h_l2213_c2_3307_cond;
     t8_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue;
     t8_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2213_c2_3307_return_output := t8_MUX_uxn_opcodes_h_l2213_c2_3307_return_output;

     -- n8_MUX[uxn_opcodes_h_l2226_c7_41d8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2226_c7_41d8_cond <= VAR_n8_MUX_uxn_opcodes_h_l2226_c7_41d8_cond;
     n8_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue;
     n8_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output := n8_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2226_c7_41d8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2233_c7_a443] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_cond;
     tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_return_output := tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2233_c7_a443] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_return_output := result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2226_c7_41d8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2226_c7_41d8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2226_c7_41d8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_a443_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2213_c2_3307_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_a443_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l2229_c7_ad46] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_cond;
     tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output := tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2229_c7_ad46] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output := result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2213_c2_3307] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2213_c2_3307] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2213_c2_3307] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2213_c2_3307] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_return_output;

     -- n8_MUX[uxn_opcodes_h_l2213_c2_3307] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2213_c2_3307_cond <= VAR_n8_MUX_uxn_opcodes_h_l2213_c2_3307_cond;
     n8_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue;
     n8_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2213_c2_3307_return_output := n8_MUX_uxn_opcodes_h_l2213_c2_3307_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2213_c2_3307_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_ad46_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2226_c7_41d8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output := result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2226_c7_41d8] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_cond;
     tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output := tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output;

     -- Submodule level 6
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_41d8_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l2213_c2_3307] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_cond;
     tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_return_output := tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2213_c2_3307] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_return_output := result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_return_output;

     -- Submodule level 7
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_3307_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l2243_l2209_DUPLICATE_685e LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l2243_l2209_DUPLICATE_685e_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6(
     result,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_3307_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_3307_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_3307_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_3307_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_3307_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_3307_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_3307_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_3307_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_3307_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l2243_l2209_DUPLICATE_685e_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l2243_l2209_DUPLICATE_685e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
