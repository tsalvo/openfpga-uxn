-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 53
entity equ_0CLK_6d7675a8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end equ_0CLK_6d7675a8;
architecture arch of equ_0CLK_6d7675a8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1231_c6_cf2f]
signal BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1231_c1_fbe1]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1231_c2_5d17]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1231_c2_5d17]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1231_c2_5d17]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1231_c2_5d17]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1231_c2_5d17]
signal result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1231_c2_5d17]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1231_c2_5d17]
signal t8_MUX_uxn_opcodes_h_l1231_c2_5d17_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1231_c2_5d17]
signal n8_MUX_uxn_opcodes_h_l1231_c2_5d17_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1232_c3_fe61[uxn_opcodes_h_l1232_c3_fe61]
signal printf_uxn_opcodes_h_l1232_c3_fe61_uxn_opcodes_h_l1232_c3_fe61_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1236_c11_eb38]
signal BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1236_c7_50f1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1236_c7_50f1]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1236_c7_50f1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1236_c7_50f1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1236_c7_50f1]
signal result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1236_c7_50f1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1236_c7_50f1]
signal t8_MUX_uxn_opcodes_h_l1236_c7_50f1_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1236_c7_50f1]
signal n8_MUX_uxn_opcodes_h_l1236_c7_50f1_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1239_c11_f1f9]
signal BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1239_c7_ee22]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1239_c7_ee22]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1239_c7_ee22]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1239_c7_ee22]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1239_c7_ee22]
signal result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1239_c7_ee22]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1239_c7_ee22]
signal t8_MUX_uxn_opcodes_h_l1239_c7_ee22_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1239_c7_ee22]
signal n8_MUX_uxn_opcodes_h_l1239_c7_ee22_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1243_c11_7135]
signal BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1243_c7_2c28]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1243_c7_2c28]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1243_c7_2c28]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1243_c7_2c28]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1243_c7_2c28]
signal result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1243_c7_2c28]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l1243_c7_2c28]
signal n8_MUX_uxn_opcodes_h_l1243_c7_2c28_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1246_c11_5b27]
signal BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1246_c7_c919]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1246_c7_c919]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1246_c7_c919]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1246_c7_c919]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1246_c7_c919]
signal result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1246_c7_c919]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l1246_c7_c919]
signal n8_MUX_uxn_opcodes_h_l1246_c7_c919_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1246_c7_c919_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1249_c30_4e8f]
signal sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1252_c21_0e0b]
signal BIN_OP_EQ_uxn_opcodes_h_l1252_c21_0e0b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1252_c21_0e0b_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1252_c21_0e0b_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1252_c21_6186]
signal MUX_uxn_opcodes_h_l1252_c21_6186_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1252_c21_6186_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1252_c21_6186_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1252_c21_6186_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1254_c11_f0ba]
signal BIN_OP_EQ_uxn_opcodes_h_l1254_c11_f0ba_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1254_c11_f0ba_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1254_c11_f0ba_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1254_c7_e719]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1254_c7_e719]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1254_c7_e719]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_641b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f
BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_left,
BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_right,
BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17
result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17
result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17
result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17
result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_cond,
result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17
result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output);

-- t8_MUX_uxn_opcodes_h_l1231_c2_5d17
t8_MUX_uxn_opcodes_h_l1231_c2_5d17 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1231_c2_5d17_cond,
t8_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue,
t8_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse,
t8_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output);

-- n8_MUX_uxn_opcodes_h_l1231_c2_5d17
n8_MUX_uxn_opcodes_h_l1231_c2_5d17 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1231_c2_5d17_cond,
n8_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue,
n8_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse,
n8_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output);

-- printf_uxn_opcodes_h_l1232_c3_fe61_uxn_opcodes_h_l1232_c3_fe61
printf_uxn_opcodes_h_l1232_c3_fe61_uxn_opcodes_h_l1232_c3_fe61 : entity work.printf_uxn_opcodes_h_l1232_c3_fe61_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1232_c3_fe61_uxn_opcodes_h_l1232_c3_fe61_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38
BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_left,
BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_right,
BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1
result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1
result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1
result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1
result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_cond,
result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1
result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output);

-- t8_MUX_uxn_opcodes_h_l1236_c7_50f1
t8_MUX_uxn_opcodes_h_l1236_c7_50f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1236_c7_50f1_cond,
t8_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue,
t8_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse,
t8_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output);

-- n8_MUX_uxn_opcodes_h_l1236_c7_50f1
n8_MUX_uxn_opcodes_h_l1236_c7_50f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1236_c7_50f1_cond,
n8_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue,
n8_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse,
n8_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9
BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_left,
BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_right,
BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22
result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22
result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22
result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22
result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_cond,
result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22
result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output);

-- t8_MUX_uxn_opcodes_h_l1239_c7_ee22
t8_MUX_uxn_opcodes_h_l1239_c7_ee22 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1239_c7_ee22_cond,
t8_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue,
t8_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse,
t8_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output);

-- n8_MUX_uxn_opcodes_h_l1239_c7_ee22
n8_MUX_uxn_opcodes_h_l1239_c7_ee22 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1239_c7_ee22_cond,
n8_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue,
n8_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse,
n8_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135
BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_left,
BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_right,
BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28
result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28
result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28
result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28
result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_cond,
result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28
result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output);

-- n8_MUX_uxn_opcodes_h_l1243_c7_2c28
n8_MUX_uxn_opcodes_h_l1243_c7_2c28 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1243_c7_2c28_cond,
n8_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue,
n8_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse,
n8_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27
BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_left,
BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_right,
BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919
result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919
result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919
result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919
result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_cond,
result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919
result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_return_output);

-- n8_MUX_uxn_opcodes_h_l1246_c7_c919
n8_MUX_uxn_opcodes_h_l1246_c7_c919 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1246_c7_c919_cond,
n8_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue,
n8_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse,
n8_MUX_uxn_opcodes_h_l1246_c7_c919_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f
sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_ins,
sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_x,
sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_y,
sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1252_c21_0e0b
BIN_OP_EQ_uxn_opcodes_h_l1252_c21_0e0b : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1252_c21_0e0b_left,
BIN_OP_EQ_uxn_opcodes_h_l1252_c21_0e0b_right,
BIN_OP_EQ_uxn_opcodes_h_l1252_c21_0e0b_return_output);

-- MUX_uxn_opcodes_h_l1252_c21_6186
MUX_uxn_opcodes_h_l1252_c21_6186 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1252_c21_6186_cond,
MUX_uxn_opcodes_h_l1252_c21_6186_iftrue,
MUX_uxn_opcodes_h_l1252_c21_6186_iffalse,
MUX_uxn_opcodes_h_l1252_c21_6186_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1254_c11_f0ba
BIN_OP_EQ_uxn_opcodes_h_l1254_c11_f0ba : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1254_c11_f0ba_left,
BIN_OP_EQ_uxn_opcodes_h_l1254_c11_f0ba_right,
BIN_OP_EQ_uxn_opcodes_h_l1254_c11_f0ba_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719
result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719
result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719
result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output,
 t8_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output,
 n8_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output,
 t8_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output,
 n8_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output,
 t8_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output,
 n8_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output,
 n8_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_return_output,
 n8_MUX_uxn_opcodes_h_l1246_c7_c919_return_output,
 sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1252_c21_0e0b_return_output,
 MUX_uxn_opcodes_h_l1252_c21_6186_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1254_c11_f0ba_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_iffalse : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1233_c3_52bd : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1231_c2_5d17_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1231_c2_5d17_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1232_c3_fe61_uxn_opcodes_h_l1232_c3_fe61_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1237_c3_2d0d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1236_c7_50f1_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1236_c7_50f1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1241_c3_b051 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1239_c7_ee22_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1239_c7_ee22_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1244_c3_d22a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1246_c7_c919_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1243_c7_2c28_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1251_c3_431a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1246_c7_c919_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1246_c7_c919_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1252_c21_6186_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1252_c21_6186_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1252_c21_6186_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1252_c21_0e0b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1252_c21_0e0b_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1252_c21_0e0b_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1252_c21_6186_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1254_c11_f0ba_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1254_c11_f0ba_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1254_c11_f0ba_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1236_l1231_l1243_l1239_l1254_DUPLICATE_47cd_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1236_l1231_l1243_l1239_l1254_DUPLICATE_f3dc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1246_l1236_l1231_l1243_l1239_DUPLICATE_015c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1246_l1236_l1231_l1243_l1239_DUPLICATE_702d_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1246_l1236_l1243_l1239_l1254_DUPLICATE_2c2c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1260_l1227_DUPLICATE_024c_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1254_c11_f0ba_right := to_unsigned(5, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1251_c3_431a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1251_c3_431a;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1233_c3_52bd := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1233_c3_52bd;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1252_c21_6186_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_MUX_uxn_opcodes_h_l1252_c21_6186_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1244_c3_d22a := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1244_c3_d22a;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1241_c3_b051 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1241_c3_b051;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1237_c3_2d0d := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1237_c3_2d0d;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_right := to_unsigned(3, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1254_c11_f0ba_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1252_c21_0e0b_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1252_c21_0e0b_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse := t8;
     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1246_c7_c919] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1246_c7_c919_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1246_c11_5b27] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_left;
     BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_return_output := BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1243_c11_7135] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_left;
     BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_return_output := BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1236_l1231_l1243_l1239_l1254_DUPLICATE_f3dc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1236_l1231_l1243_l1239_l1254_DUPLICATE_f3dc_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1236_c11_eb38] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_left;
     BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_return_output := BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1249_c30_4e8f] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_ins;
     sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_x;
     sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_return_output := sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1254_c11_f0ba] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1254_c11_f0ba_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1254_c11_f0ba_left;
     BIN_OP_EQ_uxn_opcodes_h_l1254_c11_f0ba_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1254_c11_f0ba_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1254_c11_f0ba_return_output := BIN_OP_EQ_uxn_opcodes_h_l1254_c11_f0ba_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1246_l1236_l1231_l1243_l1239_DUPLICATE_702d LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1246_l1236_l1231_l1243_l1239_DUPLICATE_702d_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1246_l1236_l1243_l1239_l1254_DUPLICATE_2c2c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1246_l1236_l1243_l1239_l1254_DUPLICATE_2c2c_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1252_c21_0e0b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1252_c21_0e0b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1252_c21_0e0b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1252_c21_0e0b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1252_c21_0e0b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1252_c21_0e0b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1252_c21_0e0b_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1246_l1236_l1231_l1243_l1239_DUPLICATE_015c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1246_l1236_l1231_l1243_l1239_DUPLICATE_015c_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1236_l1231_l1243_l1239_l1254_DUPLICATE_47cd LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1236_l1231_l1243_l1239_l1254_DUPLICATE_47cd_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1231_c6_cf2f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1239_c11_f1f9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_left;
     BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_return_output := BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1231_c2_5d17_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1231_c2_5d17_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1231_c6_cf2f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1236_c7_50f1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1236_c7_50f1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1236_c11_eb38_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1239_c7_ee22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1239_c7_ee22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1239_c11_f1f9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1243_c7_2c28_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1243_c11_7135_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1246_c7_c919_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1246_c11_5b27_return_output;
     VAR_MUX_uxn_opcodes_h_l1252_c21_6186_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1252_c21_0e0b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1254_c11_f0ba_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1254_c11_f0ba_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1254_c11_f0ba_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1246_l1236_l1231_l1243_l1239_DUPLICATE_702d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1246_l1236_l1231_l1243_l1239_DUPLICATE_702d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1246_l1236_l1231_l1243_l1239_DUPLICATE_702d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1246_l1236_l1231_l1243_l1239_DUPLICATE_702d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1246_l1236_l1231_l1243_l1239_DUPLICATE_702d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1246_l1236_l1243_l1239_l1254_DUPLICATE_2c2c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1246_l1236_l1243_l1239_l1254_DUPLICATE_2c2c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1246_l1236_l1243_l1239_l1254_DUPLICATE_2c2c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1246_l1236_l1243_l1239_l1254_DUPLICATE_2c2c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1246_l1236_l1243_l1239_l1254_DUPLICATE_2c2c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1236_l1231_l1243_l1239_l1254_DUPLICATE_47cd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1236_l1231_l1243_l1239_l1254_DUPLICATE_47cd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1236_l1231_l1243_l1239_l1254_DUPLICATE_47cd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1236_l1231_l1243_l1239_l1254_DUPLICATE_47cd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1236_l1231_l1243_l1239_l1254_DUPLICATE_47cd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1236_l1231_l1243_l1239_l1254_DUPLICATE_f3dc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1236_l1231_l1243_l1239_l1254_DUPLICATE_f3dc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1236_l1231_l1243_l1239_l1254_DUPLICATE_f3dc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1236_l1231_l1243_l1239_l1254_DUPLICATE_f3dc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1236_l1231_l1243_l1239_l1254_DUPLICATE_f3dc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1246_l1236_l1231_l1243_l1239_DUPLICATE_015c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1246_l1236_l1231_l1243_l1239_DUPLICATE_015c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1246_l1236_l1231_l1243_l1239_DUPLICATE_015c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1246_l1236_l1231_l1243_l1239_DUPLICATE_015c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1246_l1236_l1231_l1243_l1239_DUPLICATE_015c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1246_c7_c919_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1249_c30_4e8f_return_output;
     -- MUX[uxn_opcodes_h_l1252_c21_6186] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1252_c21_6186_cond <= VAR_MUX_uxn_opcodes_h_l1252_c21_6186_cond;
     MUX_uxn_opcodes_h_l1252_c21_6186_iftrue <= VAR_MUX_uxn_opcodes_h_l1252_c21_6186_iftrue;
     MUX_uxn_opcodes_h_l1252_c21_6186_iffalse <= VAR_MUX_uxn_opcodes_h_l1252_c21_6186_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1252_c21_6186_return_output := MUX_uxn_opcodes_h_l1252_c21_6186_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1246_c7_c919] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1254_c7_e719] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1246_c7_c919] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_return_output;

     -- t8_MUX[uxn_opcodes_h_l1239_c7_ee22] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1239_c7_ee22_cond <= VAR_t8_MUX_uxn_opcodes_h_l1239_c7_ee22_cond;
     t8_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue;
     t8_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output := t8_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1231_c1_fbe1] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1254_c7_e719] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_return_output;

     -- n8_MUX[uxn_opcodes_h_l1246_c7_c919] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1246_c7_c919_cond <= VAR_n8_MUX_uxn_opcodes_h_l1246_c7_c919_cond;
     n8_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue;
     n8_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1246_c7_c919_return_output := n8_MUX_uxn_opcodes_h_l1246_c7_c919_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1254_c7_e719] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue := VAR_MUX_uxn_opcodes_h_l1252_c21_6186_return_output;
     VAR_printf_uxn_opcodes_h_l1232_c3_fe61_uxn_opcodes_h_l1232_c3_fe61_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1231_c1_fbe1_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1246_c7_c919_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1254_c7_e719_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1254_c7_e719_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1254_c7_e719_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1246_c7_c919_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1246_c7_c919_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output;
     -- printf_uxn_opcodes_h_l1232_c3_fe61[uxn_opcodes_h_l1232_c3_fe61] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1232_c3_fe61_uxn_opcodes_h_l1232_c3_fe61_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1232_c3_fe61_uxn_opcodes_h_l1232_c3_fe61_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1246_c7_c919] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_return_output;

     -- n8_MUX[uxn_opcodes_h_l1243_c7_2c28] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1243_c7_2c28_cond <= VAR_n8_MUX_uxn_opcodes_h_l1243_c7_2c28_cond;
     n8_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue;
     n8_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output := n8_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1246_c7_c919] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1246_c7_c919] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_return_output := result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1243_c7_2c28] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1243_c7_2c28] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output;

     -- t8_MUX[uxn_opcodes_h_l1236_c7_50f1] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1236_c7_50f1_cond <= VAR_t8_MUX_uxn_opcodes_h_l1236_c7_50f1_cond;
     t8_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue;
     t8_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output := t8_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1246_c7_c919] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1246_c7_c919_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1246_c7_c919_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1246_c7_c919_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1246_c7_c919_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1243_c7_2c28] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1243_c7_2c28] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output := result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output;

     -- t8_MUX[uxn_opcodes_h_l1231_c2_5d17] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1231_c2_5d17_cond <= VAR_t8_MUX_uxn_opcodes_h_l1231_c2_5d17_cond;
     t8_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue;
     t8_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output := t8_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1239_c7_ee22] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1243_c7_2c28] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1239_c7_ee22] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1243_c7_2c28] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output;

     -- n8_MUX[uxn_opcodes_h_l1239_c7_ee22] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1239_c7_ee22_cond <= VAR_n8_MUX_uxn_opcodes_h_l1239_c7_ee22_cond;
     n8_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue;
     n8_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output := n8_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1243_c7_2c28_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1236_c7_50f1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1236_c7_50f1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1239_c7_ee22] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output := result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output;

     -- n8_MUX[uxn_opcodes_h_l1236_c7_50f1] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1236_c7_50f1_cond <= VAR_n8_MUX_uxn_opcodes_h_l1236_c7_50f1_cond;
     n8_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue;
     n8_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output := n8_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1239_c7_ee22] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1239_c7_ee22] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1239_c7_ee22] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1239_c7_ee22_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1231_c2_5d17] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1231_c2_5d17] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1236_c7_50f1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output := result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1236_c7_50f1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1236_c7_50f1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output;

     -- n8_MUX[uxn_opcodes_h_l1231_c2_5d17] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1231_c2_5d17_cond <= VAR_n8_MUX_uxn_opcodes_h_l1231_c2_5d17_cond;
     n8_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue;
     n8_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output := n8_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1236_c7_50f1] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1236_c7_50f1_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1231_c2_5d17] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1231_c2_5d17] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1231_c2_5d17] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output := result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1231_c2_5d17] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1260_l1227_DUPLICATE_024c LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1260_l1227_DUPLICATE_024c_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_641b(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1231_c2_5d17_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1260_l1227_DUPLICATE_024c_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1260_l1227_DUPLICATE_024c_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
