-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity equ_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end equ_0CLK_226c8821;
architecture arch of equ_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1163_c6_858b]
signal BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1163_c2_6998]
signal t8_MUX_uxn_opcodes_h_l1163_c2_6998_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1163_c2_6998_return_output : unsigned(7 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1163_c2_6998]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1163_c2_6998]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1163_c2_6998]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1163_c2_6998]
signal result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1163_c2_6998]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1163_c2_6998]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_return_output : unsigned(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1163_c2_6998]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1163_c2_6998]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1163_c2_6998]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l1163_c2_6998]
signal n8_MUX_uxn_opcodes_h_l1163_c2_6998_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1163_c2_6998_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1176_c11_fc6f]
signal BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1176_c7_80ca]
signal t8_MUX_uxn_opcodes_h_l1176_c7_80ca_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1176_c7_80ca]
signal result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1176_c7_80ca]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1176_c7_80ca]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1176_c7_80ca]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1176_c7_80ca]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l1176_c7_80ca]
signal n8_MUX_uxn_opcodes_h_l1176_c7_80ca_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1179_c11_4c00]
signal BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1179_c7_05e4]
signal t8_MUX_uxn_opcodes_h_l1179_c7_05e4_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1179_c7_05e4]
signal result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1179_c7_05e4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1179_c7_05e4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1179_c7_05e4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1179_c7_05e4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l1179_c7_05e4]
signal n8_MUX_uxn_opcodes_h_l1179_c7_05e4_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1182_c11_8933]
signal BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1182_c7_5354]
signal result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1182_c7_5354]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1182_c7_5354]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1182_c7_5354]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1182_c7_5354]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l1182_c7_5354]
signal n8_MUX_uxn_opcodes_h_l1182_c7_5354_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1182_c7_5354_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1184_c30_cb82]
signal sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1187_c21_cebe]
signal BIN_OP_EQ_uxn_opcodes_h_l1187_c21_cebe_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1187_c21_cebe_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1187_c21_cebe_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1187_c21_85b2]
signal MUX_uxn_opcodes_h_l1187_c21_85b2_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1187_c21_85b2_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1187_c21_85b2_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1187_c21_85b2_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_375c( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_vram_write := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;
      base.is_ram_write := ref_toks_7;
      base.is_stack_index_flipped := ref_toks_8;
      base.sp_relative_shift := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b
BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_left,
BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_right,
BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_return_output);

-- t8_MUX_uxn_opcodes_h_l1163_c2_6998
t8_MUX_uxn_opcodes_h_l1163_c2_6998 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1163_c2_6998_cond,
t8_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue,
t8_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse,
t8_MUX_uxn_opcodes_h_l1163_c2_6998_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998
result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998
result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998
result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998
result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_cond,
result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998
result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998
result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998
result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_return_output);

-- n8_MUX_uxn_opcodes_h_l1163_c2_6998
n8_MUX_uxn_opcodes_h_l1163_c2_6998 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1163_c2_6998_cond,
n8_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue,
n8_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse,
n8_MUX_uxn_opcodes_h_l1163_c2_6998_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f
BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_left,
BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_right,
BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_return_output);

-- t8_MUX_uxn_opcodes_h_l1176_c7_80ca
t8_MUX_uxn_opcodes_h_l1176_c7_80ca : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1176_c7_80ca_cond,
t8_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue,
t8_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse,
t8_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca
result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_cond,
result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca
result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca
result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca
result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output);

-- n8_MUX_uxn_opcodes_h_l1176_c7_80ca
n8_MUX_uxn_opcodes_h_l1176_c7_80ca : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1176_c7_80ca_cond,
n8_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue,
n8_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse,
n8_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00
BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_left,
BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_right,
BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_return_output);

-- t8_MUX_uxn_opcodes_h_l1179_c7_05e4
t8_MUX_uxn_opcodes_h_l1179_c7_05e4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1179_c7_05e4_cond,
t8_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue,
t8_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse,
t8_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4
result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_cond,
result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4
result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4
result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4
result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output);

-- n8_MUX_uxn_opcodes_h_l1179_c7_05e4
n8_MUX_uxn_opcodes_h_l1179_c7_05e4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1179_c7_05e4_cond,
n8_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue,
n8_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse,
n8_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933
BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933_left,
BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933_right,
BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354
result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_cond,
result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354
result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354
result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354
result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_return_output);

-- n8_MUX_uxn_opcodes_h_l1182_c7_5354
n8_MUX_uxn_opcodes_h_l1182_c7_5354 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1182_c7_5354_cond,
n8_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue,
n8_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse,
n8_MUX_uxn_opcodes_h_l1182_c7_5354_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82
sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_ins,
sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_x,
sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_y,
sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1187_c21_cebe
BIN_OP_EQ_uxn_opcodes_h_l1187_c21_cebe : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1187_c21_cebe_left,
BIN_OP_EQ_uxn_opcodes_h_l1187_c21_cebe_right,
BIN_OP_EQ_uxn_opcodes_h_l1187_c21_cebe_return_output);

-- MUX_uxn_opcodes_h_l1187_c21_85b2
MUX_uxn_opcodes_h_l1187_c21_85b2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1187_c21_85b2_cond,
MUX_uxn_opcodes_h_l1187_c21_85b2_iftrue,
MUX_uxn_opcodes_h_l1187_c21_85b2_iffalse,
MUX_uxn_opcodes_h_l1187_c21_85b2_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_return_output,
 t8_MUX_uxn_opcodes_h_l1163_c2_6998_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_return_output,
 n8_MUX_uxn_opcodes_h_l1163_c2_6998_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_return_output,
 t8_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output,
 n8_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_return_output,
 t8_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output,
 n8_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_return_output,
 n8_MUX_uxn_opcodes_h_l1182_c7_5354_return_output,
 sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1187_c21_cebe_return_output,
 MUX_uxn_opcodes_h_l1187_c21_85b2_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1163_c2_6998_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1163_c2_6998_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1163_c2_6998_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1163_c2_6998_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1173_c3_2c3f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1163_c2_6998_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1163_c2_6998_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1168_c3_05d8 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1163_c2_6998_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1163_c2_6998_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1176_c7_80ca_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1177_c3_e041 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1176_c7_80ca_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1179_c7_05e4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1182_c7_5354_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1179_c7_05e4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1186_c3_08b6 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1182_c7_5354_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1187_c21_85b2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_cebe_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_cebe_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_cebe_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1187_c21_85b2_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1187_c21_85b2_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1187_c21_85b2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1163_l1182_l1176_l1179_DUPLICATE_5f0c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_b995_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_d407_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_1bdc_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1182_l1179_DUPLICATE_7c17_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_375c_uxn_opcodes_h_l1191_l1159_DUPLICATE_5b25_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1173_c3_2c3f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1173_c3_2c3f;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1177_c3_e041 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1177_c3_e041;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1187_c21_85b2_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1168_c3_05d8 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1168_c3_05d8;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1186_c3_08b6 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1186_c3_08b6;
     VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1187_c21_85b2_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_cebe_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_cebe_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1176_c11_fc6f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1163_l1182_l1176_l1179_DUPLICATE_5f0c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1163_l1182_l1176_l1179_DUPLICATE_5f0c_return_output := result.u8_value;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1163_c2_6998] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1163_c2_6998_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1179_c11_4c00] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_left;
     BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_return_output := BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1182_c11_8933] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933_left;
     BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933_return_output := BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1163_c2_6998] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1163_c2_6998_return_output := result.is_pc_updated;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_1bdc LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_1bdc_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1182_l1179_DUPLICATE_7c17 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1182_l1179_DUPLICATE_7c17_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1163_c6_858b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1187_c21_cebe] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1187_c21_cebe_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_cebe_left;
     BIN_OP_EQ_uxn_opcodes_h_l1187_c21_cebe_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_cebe_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_cebe_return_output := BIN_OP_EQ_uxn_opcodes_h_l1187_c21_cebe_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_d407 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_d407_return_output := result.is_stack_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1163_c2_6998] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1163_c2_6998_return_output := result.is_stack_index_flipped;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1163_c2_6998] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1163_c2_6998_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_b995 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_b995_return_output := result.is_opc_done;

     -- sp_relative_shift[uxn_opcodes_h_l1184_c30_cb82] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_ins;
     sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_x;
     sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_return_output := sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1163_c2_6998_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1163_c2_6998_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_858b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1176_c7_80ca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1176_c7_80ca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_fc6f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1179_c7_05e4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1179_c7_05e4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_4c00_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1182_c7_5354_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_8933_return_output;
     VAR_MUX_uxn_opcodes_h_l1187_c21_85b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_cebe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_1bdc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_1bdc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_1bdc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_b995_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_b995_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_b995_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_d407_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_d407_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_d407_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1182_l1179_DUPLICATE_7c17_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1182_l1179_DUPLICATE_7c17_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1163_l1182_l1176_l1179_DUPLICATE_5f0c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1163_l1182_l1176_l1179_DUPLICATE_5f0c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1163_l1182_l1176_l1179_DUPLICATE_5f0c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1163_l1182_l1176_l1179_DUPLICATE_5f0c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1163_c2_6998_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1163_c2_6998_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1163_c2_6998_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1163_c2_6998_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_cb82_return_output;
     -- MUX[uxn_opcodes_h_l1187_c21_85b2] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1187_c21_85b2_cond <= VAR_MUX_uxn_opcodes_h_l1187_c21_85b2_cond;
     MUX_uxn_opcodes_h_l1187_c21_85b2_iftrue <= VAR_MUX_uxn_opcodes_h_l1187_c21_85b2_iftrue;
     MUX_uxn_opcodes_h_l1187_c21_85b2_iffalse <= VAR_MUX_uxn_opcodes_h_l1187_c21_85b2_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1187_c21_85b2_return_output := MUX_uxn_opcodes_h_l1187_c21_85b2_return_output;

     -- t8_MUX[uxn_opcodes_h_l1179_c7_05e4] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1179_c7_05e4_cond <= VAR_t8_MUX_uxn_opcodes_h_l1179_c7_05e4_cond;
     t8_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue;
     t8_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output := t8_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output;

     -- n8_MUX[uxn_opcodes_h_l1182_c7_5354] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1182_c7_5354_cond <= VAR_n8_MUX_uxn_opcodes_h_l1182_c7_5354_cond;
     n8_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue;
     n8_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1182_c7_5354_return_output := n8_MUX_uxn_opcodes_h_l1182_c7_5354_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1163_c2_6998] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1163_c2_6998] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1163_c2_6998] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1163_c2_6998] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1182_c7_5354] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1182_c7_5354] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1182_c7_5354] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1182_c7_5354] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue := VAR_MUX_uxn_opcodes_h_l1187_c21_85b2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1182_c7_5354_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_5354_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_5354_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_5354_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_5354_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1179_c7_05e4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1182_c7_5354] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_return_output := result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1179_c7_05e4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1179_c7_05e4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output;

     -- n8_MUX[uxn_opcodes_h_l1179_c7_05e4] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1179_c7_05e4_cond <= VAR_n8_MUX_uxn_opcodes_h_l1179_c7_05e4_cond;
     n8_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue;
     n8_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output := n8_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1179_c7_05e4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output;

     -- t8_MUX[uxn_opcodes_h_l1176_c7_80ca] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1176_c7_80ca_cond <= VAR_t8_MUX_uxn_opcodes_h_l1176_c7_80ca_cond;
     t8_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue;
     t8_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output := t8_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_5354_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1176_c7_80ca] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1176_c7_80ca] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1179_c7_05e4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output := result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1176_c7_80ca] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output;

     -- n8_MUX[uxn_opcodes_h_l1176_c7_80ca] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1176_c7_80ca_cond <= VAR_n8_MUX_uxn_opcodes_h_l1176_c7_80ca_cond;
     n8_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue;
     n8_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output := n8_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output;

     -- t8_MUX[uxn_opcodes_h_l1163_c2_6998] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1163_c2_6998_cond <= VAR_t8_MUX_uxn_opcodes_h_l1163_c2_6998_cond;
     t8_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue;
     t8_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1163_c2_6998_return_output := t8_MUX_uxn_opcodes_h_l1163_c2_6998_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1176_c7_80ca] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_05e4_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1163_c2_6998_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1176_c7_80ca] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output := result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1163_c2_6998] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1163_c2_6998] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_return_output;

     -- n8_MUX[uxn_opcodes_h_l1163_c2_6998] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1163_c2_6998_cond <= VAR_n8_MUX_uxn_opcodes_h_l1163_c2_6998_cond;
     n8_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue;
     n8_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1163_c2_6998_return_output := n8_MUX_uxn_opcodes_h_l1163_c2_6998_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1163_c2_6998] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1163_c2_6998] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1163_c2_6998_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_80ca_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1163_c2_6998] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_return_output := result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_375c_uxn_opcodes_h_l1191_l1159_DUPLICATE_5b25 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_375c_uxn_opcodes_h_l1191_l1159_DUPLICATE_5b25_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_375c(
     result,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_6998_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_6998_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_6998_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_6998_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_6998_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_6998_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_6998_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_6998_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_6998_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_375c_uxn_opcodes_h_l1191_l1159_DUPLICATE_5b25_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_375c_uxn_opcodes_h_l1191_l1159_DUPLICATE_5b25_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
