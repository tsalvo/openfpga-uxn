-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity opc_lth_phased_0CLK_2ca51e56 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(3 downto 0);
 pc : in unsigned(15 downto 0);
 sp : in unsigned(7 downto 0);
 stack_index : in unsigned(0 downto 0);
 ins : in unsigned(7 downto 0);
 k : in unsigned(7 downto 0);
 return_output : out unsigned(0 downto 0));
end opc_lth_phased_0CLK_2ca51e56;
architecture arch of opc_lth_phased_0CLK_2ca51e56 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : unsigned(0 downto 0) := to_unsigned(0, 1);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : unsigned(0 downto 0);

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_phased_h_l508_c6_6d2c]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l508_c1_9776]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l511_c7_fbaa]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l508_c2_4614]
signal t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l508_c2_4614]
signal n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l508_c2_4614]
signal result_MUX_uxn_opcodes_phased_h_l508_c2_4614_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l508_c2_4614_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l508_c2_4614_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l508_c2_4614_return_output : unsigned(0 downto 0);

-- set_will_fail[uxn_opcodes_phased_h_l509_c12_74ac]
signal set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_sp : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_k : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_mul : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_add : signed(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l511_c11_21c0]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l511_c1_a5a6]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l514_c7_7e6b]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l511_c7_fbaa]
signal t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l511_c7_fbaa]
signal n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l511_c7_fbaa]
signal result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output : unsigned(0 downto 0);

-- t_register[uxn_opcodes_phased_h_l512_c8_721b]
signal t_register_uxn_opcodes_phased_h_l512_c8_721b_CLOCK_ENABLE : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l512_c8_721b_stack_index : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l512_c8_721b_stack_ptr : unsigned(7 downto 0);
signal t_register_uxn_opcodes_phased_h_l512_c8_721b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l514_c11_1478]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l514_c1_3748]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l517_c7_92eb]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l514_c7_7e6b]
signal t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l514_c7_7e6b]
signal n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l514_c7_7e6b]
signal result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output : unsigned(0 downto 0);

-- n_register[uxn_opcodes_phased_h_l515_c8_cb9c]
signal n_register_uxn_opcodes_phased_h_l515_c8_cb9c_CLOCK_ENABLE : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l515_c8_cb9c_stack_index : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l515_c8_cb9c_stack_ptr : unsigned(7 downto 0);
signal n_register_uxn_opcodes_phased_h_l515_c8_cb9c_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l517_c11_c1f5]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l517_c11_c1f5_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l517_c11_c1f5_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l517_c11_c1f5_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l517_c1_9444]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l520_c7_46d9]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l517_c7_92eb]
signal n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l517_c7_92eb]
signal result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_return_output : unsigned(0 downto 0);

-- n_register[uxn_opcodes_phased_h_l518_c8_7084]
signal n_register_uxn_opcodes_phased_h_l518_c8_7084_CLOCK_ENABLE : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l518_c8_7084_stack_index : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l518_c8_7084_stack_ptr : unsigned(7 downto 0);
signal n_register_uxn_opcodes_phased_h_l518_c8_7084_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l520_c11_193a]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l520_c11_193a_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l520_c11_193a_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l520_c11_193a_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l520_c1_bb16]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l523_c7_30c8]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l520_c7_46d9]
signal result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_return_output : unsigned(0 downto 0);

-- set[uxn_opcodes_phased_h_l521_c3_2b82]
signal set_uxn_opcodes_phased_h_l521_c3_2b82_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l521_c3_2b82_sp : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l521_c3_2b82_stack_index : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l521_c3_2b82_ins : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l521_c3_2b82_k : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l521_c3_2b82_mul : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l521_c3_2b82_add : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l523_c11_d901]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l523_c11_d901_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l523_c11_d901_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l523_c11_d901_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l523_c1_137a]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l523_c7_30c8]
signal result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_return_output : unsigned(0 downto 0);

-- BIN_OP_LT[uxn_opcodes_phased_h_l524_c33_51ab]
signal BIN_OP_LT_uxn_opcodes_phased_h_l524_c33_51ab_left : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_phased_h_l524_c33_51ab_right : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_phased_h_l524_c33_51ab_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_phased_h_l524_c33_1b3d]
signal MUX_uxn_opcodes_phased_h_l524_c33_1b3d_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_phased_h_l524_c33_1b3d_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_phased_h_l524_c33_1b3d_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_phased_h_l524_c33_1b3d_return_output : unsigned(7 downto 0);

-- put_stack[uxn_opcodes_phased_h_l524_c3_e3f0]
signal put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_CLOCK_ENABLE : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_sp : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_stack_index : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_offset : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_value : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l526_c11_3c96]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l526_c11_3c96_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l526_c11_3c96_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l526_c11_3c96_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l526_c7_0f1c]
signal result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_return_output : unsigned(0 downto 0);


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c
BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l508_c2_4614
t8_MUX_uxn_opcodes_phased_h_l508_c2_4614 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_cond,
t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_iftrue,
t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_iffalse,
t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l508_c2_4614
n8_MUX_uxn_opcodes_phased_h_l508_c2_4614 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_cond,
n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_iftrue,
n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_iffalse,
n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_return_output);

-- result_MUX_uxn_opcodes_phased_h_l508_c2_4614
result_MUX_uxn_opcodes_phased_h_l508_c2_4614 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l508_c2_4614_cond,
result_MUX_uxn_opcodes_phased_h_l508_c2_4614_iftrue,
result_MUX_uxn_opcodes_phased_h_l508_c2_4614_iffalse,
result_MUX_uxn_opcodes_phased_h_l508_c2_4614_return_output);

-- set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac
set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac : entity work.set_will_fail_0CLK_23eb2db7 port map (
clk,
set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_CLOCK_ENABLE,
set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_sp,
set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_k,
set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_mul,
set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_add,
set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0
BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0 : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa
t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_cond,
t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iftrue,
t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iffalse,
t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa
n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_cond,
n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iftrue,
n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iffalse,
n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output);

-- result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa
result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_cond,
result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iftrue,
result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iffalse,
result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output);

-- t_register_uxn_opcodes_phased_h_l512_c8_721b
t_register_uxn_opcodes_phased_h_l512_c8_721b : entity work.t_register_0CLK_621d5f60 port map (
clk,
t_register_uxn_opcodes_phased_h_l512_c8_721b_CLOCK_ENABLE,
t_register_uxn_opcodes_phased_h_l512_c8_721b_stack_index,
t_register_uxn_opcodes_phased_h_l512_c8_721b_stack_ptr,
t_register_uxn_opcodes_phased_h_l512_c8_721b_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478
BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b
t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_cond,
t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iftrue,
t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iffalse,
t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b
n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_cond,
n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iftrue,
n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iffalse,
n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output);

-- result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b
result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_cond,
result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iftrue,
result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iffalse,
result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output);

-- n_register_uxn_opcodes_phased_h_l515_c8_cb9c
n_register_uxn_opcodes_phased_h_l515_c8_cb9c : entity work.n_register_0CLK_621d5f60 port map (
clk,
n_register_uxn_opcodes_phased_h_l515_c8_cb9c_CLOCK_ENABLE,
n_register_uxn_opcodes_phased_h_l515_c8_cb9c_stack_index,
n_register_uxn_opcodes_phased_h_l515_c8_cb9c_stack_ptr,
n_register_uxn_opcodes_phased_h_l515_c8_cb9c_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l517_c11_c1f5
BIN_OP_EQ_uxn_opcodes_phased_h_l517_c11_c1f5 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l517_c11_c1f5_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l517_c11_c1f5_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l517_c11_c1f5_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb
n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_cond,
n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iftrue,
n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iffalse,
n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_return_output);

-- result_MUX_uxn_opcodes_phased_h_l517_c7_92eb
result_MUX_uxn_opcodes_phased_h_l517_c7_92eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_cond,
result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iftrue,
result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iffalse,
result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_return_output);

-- n_register_uxn_opcodes_phased_h_l518_c8_7084
n_register_uxn_opcodes_phased_h_l518_c8_7084 : entity work.n_register_0CLK_621d5f60 port map (
clk,
n_register_uxn_opcodes_phased_h_l518_c8_7084_CLOCK_ENABLE,
n_register_uxn_opcodes_phased_h_l518_c8_7084_stack_index,
n_register_uxn_opcodes_phased_h_l518_c8_7084_stack_ptr,
n_register_uxn_opcodes_phased_h_l518_c8_7084_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l520_c11_193a
BIN_OP_EQ_uxn_opcodes_phased_h_l520_c11_193a : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l520_c11_193a_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l520_c11_193a_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l520_c11_193a_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_return_output);

-- result_MUX_uxn_opcodes_phased_h_l520_c7_46d9
result_MUX_uxn_opcodes_phased_h_l520_c7_46d9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_cond,
result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_iftrue,
result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_iffalse,
result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_return_output);

-- set_uxn_opcodes_phased_h_l521_c3_2b82
set_uxn_opcodes_phased_h_l521_c3_2b82 : entity work.set_0CLK_6f2c5aad port map (
clk,
set_uxn_opcodes_phased_h_l521_c3_2b82_CLOCK_ENABLE,
set_uxn_opcodes_phased_h_l521_c3_2b82_sp,
set_uxn_opcodes_phased_h_l521_c3_2b82_stack_index,
set_uxn_opcodes_phased_h_l521_c3_2b82_ins,
set_uxn_opcodes_phased_h_l521_c3_2b82_k,
set_uxn_opcodes_phased_h_l521_c3_2b82_mul,
set_uxn_opcodes_phased_h_l521_c3_2b82_add);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l523_c11_d901
BIN_OP_EQ_uxn_opcodes_phased_h_l523_c11_d901 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l523_c11_d901_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l523_c11_d901_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l523_c11_d901_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_return_output);

-- result_MUX_uxn_opcodes_phased_h_l523_c7_30c8
result_MUX_uxn_opcodes_phased_h_l523_c7_30c8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_cond,
result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_iftrue,
result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_iffalse,
result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_return_output);

-- BIN_OP_LT_uxn_opcodes_phased_h_l524_c33_51ab
BIN_OP_LT_uxn_opcodes_phased_h_l524_c33_51ab : entity work.BIN_OP_LT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_LT_uxn_opcodes_phased_h_l524_c33_51ab_left,
BIN_OP_LT_uxn_opcodes_phased_h_l524_c33_51ab_right,
BIN_OP_LT_uxn_opcodes_phased_h_l524_c33_51ab_return_output);

-- MUX_uxn_opcodes_phased_h_l524_c33_1b3d
MUX_uxn_opcodes_phased_h_l524_c33_1b3d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_phased_h_l524_c33_1b3d_cond,
MUX_uxn_opcodes_phased_h_l524_c33_1b3d_iftrue,
MUX_uxn_opcodes_phased_h_l524_c33_1b3d_iffalse,
MUX_uxn_opcodes_phased_h_l524_c33_1b3d_return_output);

-- put_stack_uxn_opcodes_phased_h_l524_c3_e3f0
put_stack_uxn_opcodes_phased_h_l524_c3_e3f0 : entity work.put_stack_0CLK_b888155f port map (
clk,
put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_CLOCK_ENABLE,
put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_sp,
put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_stack_index,
put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_offset,
put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_value);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l526_c11_3c96
BIN_OP_EQ_uxn_opcodes_phased_h_l526_c11_3c96 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l526_c11_3c96_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l526_c11_3c96_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l526_c11_3c96_return_output);

-- result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c
result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_cond,
result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_iftrue,
result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_iffalse,
result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 sp,
 stack_index,
 ins,
 k,
 -- Registers
 n8,
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output,
 t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_return_output,
 n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_return_output,
 result_MUX_uxn_opcodes_phased_h_l508_c2_4614_return_output,
 set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output,
 t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output,
 n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output,
 result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output,
 t_register_uxn_opcodes_phased_h_l512_c8_721b_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_return_output,
 t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output,
 n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output,
 result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output,
 n_register_uxn_opcodes_phased_h_l515_c8_cb9c_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l517_c11_c1f5_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_return_output,
 n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_return_output,
 result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_return_output,
 n_register_uxn_opcodes_phased_h_l518_c8_7084_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l520_c11_193a_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_return_output,
 result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l523_c11_d901_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_return_output,
 result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_return_output,
 BIN_OP_LT_uxn_opcodes_phased_h_l524_c33_51ab_return_output,
 MUX_uxn_opcodes_phased_h_l524_c33_1b3d_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l526_c11_3c96_return_output,
 result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(0 downto 0);
 variable VAR_phase : unsigned(3 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_sp : unsigned(7 downto 0);
 variable VAR_stack_index : unsigned(0 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_k : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l508_c2_4614_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l508_c2_4614_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l508_c2_4614_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l508_c2_4614_cond : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_sp : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_k : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_mul : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_add : signed(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_cond : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l512_c8_721b_stack_index : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l512_c8_721b_stack_ptr : unsigned(7 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l512_c8_721b_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l512_c8_721b_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_cond : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l515_c8_cb9c_stack_index : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l515_c8_cb9c_stack_ptr : unsigned(7 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l515_c8_cb9c_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l515_c8_cb9c_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l517_c11_c1f5_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l517_c11_c1f5_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l517_c11_c1f5_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_cond : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l518_c8_7084_stack_index : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l518_c8_7084_stack_ptr : unsigned(7 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l518_c8_7084_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l518_c8_7084_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l520_c11_193a_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l520_c11_193a_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l520_c11_193a_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_cond : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l521_c3_2b82_sp : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l521_c3_2b82_stack_index : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l521_c3_2b82_ins : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l521_c3_2b82_k : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l521_c3_2b82_mul : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l521_c3_2b82_add : signed(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l521_c3_2b82_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l523_c11_d901_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l523_c11_d901_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l523_c11_d901_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_cond : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_sp : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_stack_index : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_offset : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_value : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_phased_h_l524_c33_1b3d_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_phased_h_l524_c33_1b3d_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_phased_h_l524_c33_1b3d_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_phased_h_l524_c33_51ab_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_phased_h_l524_c33_51ab_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_phased_h_l524_c33_51ab_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_phased_h_l524_c33_1b3d_return_output : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l526_c11_3c96_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l526_c11_3c96_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l526_c11_3c96_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_cond : unsigned(0 downto 0);
 -- State registers comb logic variables
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : unsigned(0 downto 0);
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_n8 := n8;
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_iffalse := to_unsigned(0, 1);
     VAR_set_uxn_opcodes_phased_h_l521_c3_2b82_mul := resize(to_unsigned(2, 2), 8);
     VAR_MUX_uxn_opcodes_phased_h_l524_c33_1b3d_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_mul := resize(to_unsigned(2, 2), 8);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l523_c11_d901_right := to_unsigned(5, 3);
     VAR_put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_offset := resize(to_unsigned(0, 1), 8);
     VAR_MUX_uxn_opcodes_phased_h_l524_c33_1b3d_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0_right := to_unsigned(1, 1);
     VAR_set_uxn_opcodes_phased_h_l521_c3_2b82_add := resize(to_signed(-1, 2), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c_right := to_unsigned(0, 1);
     VAR_set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_add := resize(to_signed(-1, 2), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l517_c11_c1f5_right := to_unsigned(3, 2);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l526_c11_3c96_right := to_unsigned(6, 3);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iftrue := to_unsigned(0, 1);
     VAR_result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l520_c11_193a_right := to_unsigned(4, 3);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_sp := sp;
     VAR_stack_index := stack_index;
     VAR_ins := ins;
     VAR_k := k;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iffalse := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_iftrue := VAR_CLOCK_ENABLE;
     VAR_set_uxn_opcodes_phased_h_l521_c3_2b82_ins := VAR_ins;
     VAR_set_uxn_opcodes_phased_h_l521_c3_2b82_k := VAR_k;
     VAR_set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_k := VAR_k;
     VAR_BIN_OP_LT_uxn_opcodes_phased_h_l524_c33_51ab_left := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l517_c11_c1f5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l520_c11_193a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l523_c11_d901_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l526_c11_3c96_left := VAR_phase;
     VAR_result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_iffalse := result;
     VAR_n_register_uxn_opcodes_phased_h_l515_c8_cb9c_stack_ptr := VAR_sp;
     VAR_n_register_uxn_opcodes_phased_h_l518_c8_7084_stack_ptr := VAR_sp;
     VAR_put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_sp := VAR_sp;
     VAR_set_uxn_opcodes_phased_h_l521_c3_2b82_sp := VAR_sp;
     VAR_set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_sp := VAR_sp;
     VAR_t_register_uxn_opcodes_phased_h_l512_c8_721b_stack_ptr := VAR_sp;
     VAR_n_register_uxn_opcodes_phased_h_l515_c8_cb9c_stack_index := VAR_stack_index;
     VAR_n_register_uxn_opcodes_phased_h_l518_c8_7084_stack_index := VAR_stack_index;
     VAR_put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_stack_index := VAR_stack_index;
     VAR_set_uxn_opcodes_phased_h_l521_c3_2b82_stack_index := VAR_stack_index;
     VAR_t_register_uxn_opcodes_phased_h_l512_c8_721b_stack_index := VAR_stack_index;
     VAR_BIN_OP_LT_uxn_opcodes_phased_h_l524_c33_51ab_right := t8;
     VAR_t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iffalse := t8;
     -- BIN_OP_LT[uxn_opcodes_phased_h_l524_c33_51ab] LATENCY=0
     -- Inputs
     BIN_OP_LT_uxn_opcodes_phased_h_l524_c33_51ab_left <= VAR_BIN_OP_LT_uxn_opcodes_phased_h_l524_c33_51ab_left;
     BIN_OP_LT_uxn_opcodes_phased_h_l524_c33_51ab_right <= VAR_BIN_OP_LT_uxn_opcodes_phased_h_l524_c33_51ab_right;
     -- Outputs
     VAR_BIN_OP_LT_uxn_opcodes_phased_h_l524_c33_51ab_return_output := BIN_OP_LT_uxn_opcodes_phased_h_l524_c33_51ab_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l523_c11_d901] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l523_c11_d901_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l523_c11_d901_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l523_c11_d901_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l523_c11_d901_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l523_c11_d901_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l523_c11_d901_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l517_c11_c1f5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l517_c11_c1f5_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l517_c11_c1f5_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l517_c11_c1f5_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l517_c11_c1f5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l517_c11_c1f5_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l517_c11_c1f5_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l514_c11_1478] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l508_c6_6d2c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l526_c11_3c96] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l526_c11_3c96_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l526_c11_3c96_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l526_c11_3c96_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l526_c11_3c96_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l526_c11_3c96_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l526_c11_3c96_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l520_c11_193a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l520_c11_193a_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l520_c11_193a_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l520_c11_193a_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l520_c11_193a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l520_c11_193a_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l520_c11_193a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l511_c11_21c0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0_return_output;

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l508_c2_4614_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l508_c6_6d2c_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l511_c11_21c0_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l514_c11_1478_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l517_c11_c1f5_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l517_c11_c1f5_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l517_c11_c1f5_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l517_c11_c1f5_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l520_c11_193a_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l520_c11_193a_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l520_c11_193a_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l523_c11_d901_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l523_c11_d901_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l526_c11_3c96_return_output;
     VAR_MUX_uxn_opcodes_phased_h_l524_c33_1b3d_cond := VAR_BIN_OP_LT_uxn_opcodes_phased_h_l524_c33_51ab_return_output;
     -- MUX[uxn_opcodes_phased_h_l524_c33_1b3d] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_phased_h_l524_c33_1b3d_cond <= VAR_MUX_uxn_opcodes_phased_h_l524_c33_1b3d_cond;
     MUX_uxn_opcodes_phased_h_l524_c33_1b3d_iftrue <= VAR_MUX_uxn_opcodes_phased_h_l524_c33_1b3d_iftrue;
     MUX_uxn_opcodes_phased_h_l524_c33_1b3d_iffalse <= VAR_MUX_uxn_opcodes_phased_h_l524_c33_1b3d_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_phased_h_l524_c33_1b3d_return_output := MUX_uxn_opcodes_phased_h_l524_c33_1b3d_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l526_c7_0f1c] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_cond;
     result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_iftrue;
     result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_return_output := result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l511_c7_fbaa] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l508_c1_9776] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output;
     VAR_put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_value := VAR_MUX_uxn_opcodes_phased_h_l524_c33_1b3d_return_output;
     VAR_set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l508_c1_9776_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l526_c7_0f1c_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l523_c7_30c8] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_cond;
     result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_iftrue;
     result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_return_output := result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l511_c1_a5a6] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l514_c7_7e6b] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output;

     -- set_will_fail[uxn_opcodes_phased_h_l509_c12_74ac] LATENCY=0
     -- Clock enable
     set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_CLOCK_ENABLE <= VAR_set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_CLOCK_ENABLE;
     -- Inputs
     set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_sp <= VAR_set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_sp;
     set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_k <= VAR_set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_k;
     set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_mul <= VAR_set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_mul;
     set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_add <= VAR_set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_add;
     -- Outputs
     VAR_set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_return_output := set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_return_output;

     -- Submodule level 3
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output;
     VAR_t_register_uxn_opcodes_phased_h_l512_c8_721b_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l511_c1_a5a6_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l523_c7_30c8_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l508_c2_4614_iftrue := VAR_set_will_fail_uxn_opcodes_phased_h_l509_c12_74ac_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l514_c1_3748] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_return_output;

     -- t_register[uxn_opcodes_phased_h_l512_c8_721b] LATENCY=0
     -- Clock enable
     t_register_uxn_opcodes_phased_h_l512_c8_721b_CLOCK_ENABLE <= VAR_t_register_uxn_opcodes_phased_h_l512_c8_721b_CLOCK_ENABLE;
     -- Inputs
     t_register_uxn_opcodes_phased_h_l512_c8_721b_stack_index <= VAR_t_register_uxn_opcodes_phased_h_l512_c8_721b_stack_index;
     t_register_uxn_opcodes_phased_h_l512_c8_721b_stack_ptr <= VAR_t_register_uxn_opcodes_phased_h_l512_c8_721b_stack_ptr;
     -- Outputs
     VAR_t_register_uxn_opcodes_phased_h_l512_c8_721b_return_output := t_register_uxn_opcodes_phased_h_l512_c8_721b_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l520_c7_46d9] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_cond;
     result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_iftrue;
     result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_return_output := result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l517_c7_92eb] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_return_output;

     -- Submodule level 4
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c7_92eb_return_output;
     VAR_n_register_uxn_opcodes_phased_h_l515_c8_cb9c_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l514_c1_3748_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l520_c7_46d9_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iftrue := VAR_t_register_uxn_opcodes_phased_h_l512_c8_721b_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l520_c7_46d9] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l517_c1_9444] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_return_output;

     -- n_register[uxn_opcodes_phased_h_l515_c8_cb9c] LATENCY=0
     -- Clock enable
     n_register_uxn_opcodes_phased_h_l515_c8_cb9c_CLOCK_ENABLE <= VAR_n_register_uxn_opcodes_phased_h_l515_c8_cb9c_CLOCK_ENABLE;
     -- Inputs
     n_register_uxn_opcodes_phased_h_l515_c8_cb9c_stack_index <= VAR_n_register_uxn_opcodes_phased_h_l515_c8_cb9c_stack_index;
     n_register_uxn_opcodes_phased_h_l515_c8_cb9c_stack_ptr <= VAR_n_register_uxn_opcodes_phased_h_l515_c8_cb9c_stack_ptr;
     -- Outputs
     VAR_n_register_uxn_opcodes_phased_h_l515_c8_cb9c_return_output := n_register_uxn_opcodes_phased_h_l515_c8_cb9c_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l517_c7_92eb] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_cond;
     result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iftrue;
     result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_return_output := result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_return_output;

     -- Submodule level 5
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c7_46d9_return_output;
     VAR_n_register_uxn_opcodes_phased_h_l518_c8_7084_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l517_c1_9444_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iftrue := VAR_n_register_uxn_opcodes_phased_h_l515_c8_cb9c_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l517_c7_92eb_return_output;
     -- t8_MUX[uxn_opcodes_phased_h_l514_c7_7e6b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_cond;
     t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output := t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output;

     -- n_register[uxn_opcodes_phased_h_l518_c8_7084] LATENCY=0
     -- Clock enable
     n_register_uxn_opcodes_phased_h_l518_c8_7084_CLOCK_ENABLE <= VAR_n_register_uxn_opcodes_phased_h_l518_c8_7084_CLOCK_ENABLE;
     -- Inputs
     n_register_uxn_opcodes_phased_h_l518_c8_7084_stack_index <= VAR_n_register_uxn_opcodes_phased_h_l518_c8_7084_stack_index;
     n_register_uxn_opcodes_phased_h_l518_c8_7084_stack_ptr <= VAR_n_register_uxn_opcodes_phased_h_l518_c8_7084_stack_ptr;
     -- Outputs
     VAR_n_register_uxn_opcodes_phased_h_l518_c8_7084_return_output := n_register_uxn_opcodes_phased_h_l518_c8_7084_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l520_c1_bb16] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l514_c7_7e6b] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_cond;
     result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iftrue;
     result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output := result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l523_c7_30c8] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_return_output;

     -- Submodule level 6
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c7_30c8_return_output;
     VAR_set_uxn_opcodes_phased_h_l521_c3_2b82_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l520_c1_bb16_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iftrue := VAR_n_register_uxn_opcodes_phased_h_l518_c8_7084_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iffalse := VAR_t8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l523_c1_137a] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l511_c7_fbaa] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_cond;
     result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iftrue;
     result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output := result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output;

     -- t8_MUX[uxn_opcodes_phased_h_l511_c7_fbaa] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_cond;
     t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output := t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output;

     -- n8_MUX[uxn_opcodes_phased_h_l517_c7_92eb] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_cond;
     n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_return_output := n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_return_output;

     -- set[uxn_opcodes_phased_h_l521_c3_2b82] LATENCY=0
     -- Clock enable
     set_uxn_opcodes_phased_h_l521_c3_2b82_CLOCK_ENABLE <= VAR_set_uxn_opcodes_phased_h_l521_c3_2b82_CLOCK_ENABLE;
     -- Inputs
     set_uxn_opcodes_phased_h_l521_c3_2b82_sp <= VAR_set_uxn_opcodes_phased_h_l521_c3_2b82_sp;
     set_uxn_opcodes_phased_h_l521_c3_2b82_stack_index <= VAR_set_uxn_opcodes_phased_h_l521_c3_2b82_stack_index;
     set_uxn_opcodes_phased_h_l521_c3_2b82_ins <= VAR_set_uxn_opcodes_phased_h_l521_c3_2b82_ins;
     set_uxn_opcodes_phased_h_l521_c3_2b82_k <= VAR_set_uxn_opcodes_phased_h_l521_c3_2b82_k;
     set_uxn_opcodes_phased_h_l521_c3_2b82_mul <= VAR_set_uxn_opcodes_phased_h_l521_c3_2b82_mul;
     set_uxn_opcodes_phased_h_l521_c3_2b82_add <= VAR_set_uxn_opcodes_phased_h_l521_c3_2b82_add;
     -- Outputs

     -- Submodule level 7
     VAR_put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l523_c1_137a_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l517_c7_92eb_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l508_c2_4614_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_iffalse := VAR_t8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output;
     -- t8_MUX[uxn_opcodes_phased_h_l508_c2_4614] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_cond;
     t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_return_output := t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_return_output;

     -- put_stack[uxn_opcodes_phased_h_l524_c3_e3f0] LATENCY=0
     -- Clock enable
     put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_CLOCK_ENABLE <= VAR_put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_CLOCK_ENABLE;
     -- Inputs
     put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_sp <= VAR_put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_sp;
     put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_stack_index <= VAR_put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_stack_index;
     put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_offset <= VAR_put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_offset;
     put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_value <= VAR_put_stack_uxn_opcodes_phased_h_l524_c3_e3f0_value;
     -- Outputs

     -- n8_MUX[uxn_opcodes_phased_h_l514_c7_7e6b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_cond;
     n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output := n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l508_c2_4614] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l508_c2_4614_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l508_c2_4614_cond;
     result_MUX_uxn_opcodes_phased_h_l508_c2_4614_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l508_c2_4614_iftrue;
     result_MUX_uxn_opcodes_phased_h_l508_c2_4614_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l508_c2_4614_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l508_c2_4614_return_output := result_MUX_uxn_opcodes_phased_h_l508_c2_4614_return_output;

     -- Submodule level 8
     VAR_n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l514_c7_7e6b_return_output;
     REG_VAR_result := VAR_result_MUX_uxn_opcodes_phased_h_l508_c2_4614_return_output;
     VAR_return_output := VAR_result_MUX_uxn_opcodes_phased_h_l508_c2_4614_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_phased_h_l508_c2_4614_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l511_c7_fbaa] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_cond;
     n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output := n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output;

     -- Submodule level 9
     VAR_n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l511_c7_fbaa_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l508_c2_4614] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_cond;
     n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_return_output := n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_return_output;

     -- Submodule level 10
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_phased_h_l508_c2_4614_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     n8 <= REG_COMB_n8;
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
